
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY wav_rom IS
PORT (
      CLOCK          : IN  STD_LOGIC;
      ce : in std_logic;
      ADDR_1         : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
      ADDR_2 : in std_logic_vector(15 downto 0);
      two_notes : in std_logic;
      DATA_OUT       : OUT STD_LOGIC_VECTOR(10 DOWNTO 0)
      );
END wav_rom;

ARCHITECTURE Behavioral OF wav_rom IS

  TYPE rom_type IS ARRAY (0 TO 41894) OF SIGNED (10 DOWNTO 0);
  SIGNAL memory : rom_type := (
TO_SIGNED(0,11),
TO_SIGNED(47,11),
TO_SIGNED(94,11),
TO_SIGNED(140,11),
TO_SIGNED(186,11),
TO_SIGNED(231,11),
TO_SIGNED(275,11),
TO_SIGNED(319,11),
TO_SIGNED(361,11),
TO_SIGNED(401,11),
TO_SIGNED(440,11),
TO_SIGNED(477,11),
TO_SIGNED(512,11),
TO_SIGNED(546,11),
TO_SIGNED(577,11),
TO_SIGNED(606,11),
TO_SIGNED(632,11),
TO_SIGNED(656,11),
TO_SIGNED(678,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(736,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(699,11),
TO_SIGNED(680,11),
TO_SIGNED(659,11),
TO_SIGNED(635,11),
TO_SIGNED(609,11),
TO_SIGNED(580,11),
TO_SIGNED(549,11),
TO_SIGNED(516,11),
TO_SIGNED(481,11),
TO_SIGNED(444,11),
TO_SIGNED(406,11),
TO_SIGNED(365,11),
TO_SIGNED(323,11),
TO_SIGNED(280,11),
TO_SIGNED(236,11),
TO_SIGNED(191,11),
TO_SIGNED(145,11),
TO_SIGNED(99,11),
TO_SIGNED(52,11),
TO_SIGNED(5,11),
TO_SIGNED(-42,11),
TO_SIGNED(-88,11),
TO_SIGNED(-135,11),
TO_SIGNED(-181,11),
TO_SIGNED(-226,11),
TO_SIGNED(-271,11),
TO_SIGNED(-314,11),
TO_SIGNED(-356,11),
TO_SIGNED(-397,11),
TO_SIGNED(-436,11),
TO_SIGNED(-473,11),
TO_SIGNED(-509,11),
TO_SIGNED(-542,11),
TO_SIGNED(-574,11),
TO_SIGNED(-603,11),
TO_SIGNED(-629,11),
TO_SIGNED(-654,11),
TO_SIGNED(-675,11),
TO_SIGNED(-695,11),
TO_SIGNED(-711,11),
TO_SIGNED(-725,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-716,11),
TO_SIGNED(-700,11),
TO_SIGNED(-682,11),
TO_SIGNED(-661,11),
TO_SIGNED(-638,11),
TO_SIGNED(-612,11),
TO_SIGNED(-584,11),
TO_SIGNED(-553,11),
TO_SIGNED(-520,11),
TO_SIGNED(-485,11),
TO_SIGNED(-449,11),
TO_SIGNED(-410,11),
TO_SIGNED(-370,11),
TO_SIGNED(-328,11),
TO_SIGNED(-285,11),
TO_SIGNED(-241,11),
TO_SIGNED(-196,11),
TO_SIGNED(-151,11),
TO_SIGNED(-104,11),
TO_SIGNED(-58,11),
TO_SIGNED(-11,11),
TO_SIGNED(36,11),
TO_SIGNED(83,11),
TO_SIGNED(130,11),
TO_SIGNED(176,11),
TO_SIGNED(221,11),
TO_SIGNED(266,11),
TO_SIGNED(309,11),
TO_SIGNED(351,11),
TO_SIGNED(392,11),
TO_SIGNED(431,11),
TO_SIGNED(469,11),
TO_SIGNED(505,11),
TO_SIGNED(538,11),
TO_SIGNED(570,11),
TO_SIGNED(599,11),
TO_SIGNED(627,11),
TO_SIGNED(651,11),
TO_SIGNED(673,11),
TO_SIGNED(693,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(739,11),
TO_SIGNED(730,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(685,11),
TO_SIGNED(664,11),
TO_SIGNED(641,11),
TO_SIGNED(615,11),
TO_SIGNED(587,11),
TO_SIGNED(557,11),
TO_SIGNED(524,11),
TO_SIGNED(489,11),
TO_SIGNED(453,11),
TO_SIGNED(415,11),
TO_SIGNED(375,11),
TO_SIGNED(333,11),
TO_SIGNED(290,11),
TO_SIGNED(246,11),
TO_SIGNED(202,11),
TO_SIGNED(156,11),
TO_SIGNED(110,11),
TO_SIGNED(63,11),
TO_SIGNED(16,11),
TO_SIGNED(-31,11),
TO_SIGNED(-78,11),
TO_SIGNED(-124,11),
TO_SIGNED(-171,11),
TO_SIGNED(-216,11),
TO_SIGNED(-261,11),
TO_SIGNED(-304,11),
TO_SIGNED(-346,11),
TO_SIGNED(-387,11),
TO_SIGNED(-427,11),
TO_SIGNED(-465,11),
TO_SIGNED(-501,11),
TO_SIGNED(-535,11),
TO_SIGNED(-567,11),
TO_SIGNED(-596,11),
TO_SIGNED(-624,11),
TO_SIGNED(-648,11),
TO_SIGNED(-671,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-719,11),
TO_SIGNED(-704,11),
TO_SIGNED(-687,11),
TO_SIGNED(-666,11),
TO_SIGNED(-644,11),
TO_SIGNED(-618,11),
TO_SIGNED(-590,11),
TO_SIGNED(-560,11),
TO_SIGNED(-528,11),
TO_SIGNED(-493,11),
TO_SIGNED(-457,11),
TO_SIGNED(-419,11),
TO_SIGNED(-379,11),
TO_SIGNED(-338,11),
TO_SIGNED(-295,11),
TO_SIGNED(-251,11),
TO_SIGNED(-207,11),
TO_SIGNED(-161,11),
TO_SIGNED(-115,11),
TO_SIGNED(-68,11),
TO_SIGNED(-21,11),
TO_SIGNED(26,11),
TO_SIGNED(73,11),
TO_SIGNED(119,11),
TO_SIGNED(165,11),
TO_SIGNED(211,11),
TO_SIGNED(256,11),
TO_SIGNED(299,11),
TO_SIGNED(342,11),
TO_SIGNED(383,11),
TO_SIGNED(422,11),
TO_SIGNED(460,11),
TO_SIGNED(497,11),
TO_SIGNED(531,11),
TO_SIGNED(563,11),
TO_SIGNED(593,11),
TO_SIGNED(621,11),
TO_SIGNED(646,11),
TO_SIGNED(668,11),
TO_SIGNED(688,11),
TO_SIGNED(706,11),
TO_SIGNED(720,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(721,11),
TO_SIGNED(706,11),
TO_SIGNED(689,11),
TO_SIGNED(669,11),
TO_SIGNED(646,11),
TO_SIGNED(621,11),
TO_SIGNED(594,11),
TO_SIGNED(564,11),
TO_SIGNED(532,11),
TO_SIGNED(497,11),
TO_SIGNED(461,11),
TO_SIGNED(423,11),
TO_SIGNED(384,11),
TO_SIGNED(343,11),
TO_SIGNED(300,11),
TO_SIGNED(257,11),
TO_SIGNED(212,11),
TO_SIGNED(166,11),
TO_SIGNED(120,11),
TO_SIGNED(74,11),
TO_SIGNED(27,11),
TO_SIGNED(-20,11),
TO_SIGNED(-67,11),
TO_SIGNED(-114,11),
TO_SIGNED(-160,11),
TO_SIGNED(-206,11),
TO_SIGNED(-250,11),
TO_SIGNED(-294,11),
TO_SIGNED(-337,11),
TO_SIGNED(-378,11),
TO_SIGNED(-418,11),
TO_SIGNED(-456,11),
TO_SIGNED(-493,11),
TO_SIGNED(-527,11),
TO_SIGNED(-559,11),
TO_SIGNED(-590,11),
TO_SIGNED(-618,11),
TO_SIGNED(-643,11),
TO_SIGNED(-666,11),
TO_SIGNED(-686,11),
TO_SIGNED(-704,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-733,11),
TO_SIGNED(-722,11),
TO_SIGNED(-708,11),
TO_SIGNED(-691,11),
TO_SIGNED(-671,11),
TO_SIGNED(-649,11),
TO_SIGNED(-624,11),
TO_SIGNED(-597,11),
TO_SIGNED(-567,11),
TO_SIGNED(-535,11),
TO_SIGNED(-501,11),
TO_SIGNED(-466,11),
TO_SIGNED(-428,11),
TO_SIGNED(-388,11),
TO_SIGNED(-347,11),
TO_SIGNED(-305,11),
TO_SIGNED(-262,11),
TO_SIGNED(-217,11),
TO_SIGNED(-172,11),
TO_SIGNED(-125,11),
TO_SIGNED(-79,11),
TO_SIGNED(-32,11),
TO_SIGNED(15,11),
TO_SIGNED(62,11),
TO_SIGNED(109,11),
TO_SIGNED(155,11),
TO_SIGNED(201,11),
TO_SIGNED(245,11),
TO_SIGNED(289,11),
TO_SIGNED(332,11),
TO_SIGNED(374,11),
TO_SIGNED(414,11),
TO_SIGNED(452,11),
TO_SIGNED(489,11),
TO_SIGNED(523,11),
TO_SIGNED(556,11),
TO_SIGNED(586,11),
TO_SIGNED(615,11),
TO_SIGNED(640,11),
TO_SIGNED(663,11),
TO_SIGNED(684,11),
TO_SIGNED(702,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(710,11),
TO_SIGNED(693,11),
TO_SIGNED(674,11),
TO_SIGNED(652,11),
TO_SIGNED(627,11),
TO_SIGNED(600,11),
TO_SIGNED(571,11),
TO_SIGNED(539,11),
TO_SIGNED(505,11),
TO_SIGNED(470,11),
TO_SIGNED(432,11),
TO_SIGNED(393,11),
TO_SIGNED(352,11),
TO_SIGNED(310,11),
TO_SIGNED(267,11),
TO_SIGNED(222,11),
TO_SIGNED(177,11),
TO_SIGNED(131,11),
TO_SIGNED(84,11),
TO_SIGNED(37,11),
TO_SIGNED(-10,11),
TO_SIGNED(-57,11),
TO_SIGNED(-103,11),
TO_SIGNED(-150,11),
TO_SIGNED(-195,11),
TO_SIGNED(-240,11),
TO_SIGNED(-284,11),
TO_SIGNED(-327,11),
TO_SIGNED(-369,11),
TO_SIGNED(-409,11),
TO_SIGNED(-448,11),
TO_SIGNED(-485,11),
TO_SIGNED(-519,11),
TO_SIGNED(-552,11),
TO_SIGNED(-583,11),
TO_SIGNED(-611,11),
TO_SIGNED(-637,11),
TO_SIGNED(-661,11),
TO_SIGNED(-682,11),
TO_SIGNED(-700,11),
TO_SIGNED(-716,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-725,11),
TO_SIGNED(-711,11),
TO_SIGNED(-695,11),
TO_SIGNED(-676,11),
TO_SIGNED(-654,11),
TO_SIGNED(-630,11),
TO_SIGNED(-603,11),
TO_SIGNED(-574,11),
TO_SIGNED(-543,11),
TO_SIGNED(-509,11),
TO_SIGNED(-474,11),
TO_SIGNED(-437,11),
TO_SIGNED(-397,11),
TO_SIGNED(-357,11),
TO_SIGNED(-315,11),
TO_SIGNED(-272,11),
TO_SIGNED(-227,11),
TO_SIGNED(-182,11),
TO_SIGNED(-136,11),
TO_SIGNED(-90,11),
TO_SIGNED(-43,11),
TO_SIGNED(4,11),
TO_SIGNED(51,11),
TO_SIGNED(98,11),
TO_SIGNED(144,11),
TO_SIGNED(190,11),
TO_SIGNED(235,11),
TO_SIGNED(279,11),
TO_SIGNED(323,11),
TO_SIGNED(364,11),
TO_SIGNED(405,11),
TO_SIGNED(443,11),
TO_SIGNED(480,11),
TO_SIGNED(516,11),
TO_SIGNED(549,11),
TO_SIGNED(580,11),
TO_SIGNED(608,11),
TO_SIGNED(635,11),
TO_SIGNED(658,11),
TO_SIGNED(680,11),
TO_SIGNED(698,11),
TO_SIGNED(714,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(713,11),
TO_SIGNED(697,11),
TO_SIGNED(678,11),
TO_SIGNED(657,11),
TO_SIGNED(633,11),
TO_SIGNED(606,11),
TO_SIGNED(578,11),
TO_SIGNED(547,11),
TO_SIGNED(513,11),
TO_SIGNED(478,11),
TO_SIGNED(441,11),
TO_SIGNED(402,11),
TO_SIGNED(362,11),
TO_SIGNED(320,11),
TO_SIGNED(276,11),
TO_SIGNED(232,11),
TO_SIGNED(187,11),
TO_SIGNED(141,11),
TO_SIGNED(95,11),
TO_SIGNED(48,11),
TO_SIGNED(1,11),
TO_SIGNED(-46,11),
TO_SIGNED(-93,11),
TO_SIGNED(-139,11),
TO_SIGNED(-185,11),
TO_SIGNED(-230,11),
TO_SIGNED(-275,11),
TO_SIGNED(-318,11),
TO_SIGNED(-360,11),
TO_SIGNED(-400,11),
TO_SIGNED(-439,11),
TO_SIGNED(-476,11),
TO_SIGNED(-512,11),
TO_SIGNED(-545,11),
TO_SIGNED(-576,11),
TO_SIGNED(-605,11),
TO_SIGNED(-632,11),
TO_SIGNED(-656,11),
TO_SIGNED(-677,11),
TO_SIGNED(-696,11),
TO_SIGNED(-712,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-715,11),
TO_SIGNED(-699,11),
TO_SIGNED(-681,11),
TO_SIGNED(-659,11),
TO_SIGNED(-636,11),
TO_SIGNED(-610,11),
TO_SIGNED(-581,11),
TO_SIGNED(-550,11),
TO_SIGNED(-517,11),
TO_SIGNED(-482,11),
TO_SIGNED(-445,11),
TO_SIGNED(-406,11),
TO_SIGNED(-366,11),
TO_SIGNED(-324,11),
TO_SIGNED(-281,11),
TO_SIGNED(-237,11),
TO_SIGNED(-192,11),
TO_SIGNED(-147,11),
TO_SIGNED(-100,11),
TO_SIGNED(-53,11),
TO_SIGNED(-6,11),
TO_SIGNED(41,11),
TO_SIGNED(87,11),
TO_SIGNED(134,11),
TO_SIGNED(180,11),
TO_SIGNED(225,11),
TO_SIGNED(270,11),
TO_SIGNED(313,11),
TO_SIGNED(355,11),
TO_SIGNED(396,11),
TO_SIGNED(435,11),
TO_SIGNED(472,11),
TO_SIGNED(508,11),
TO_SIGNED(541,11),
TO_SIGNED(573,11),
TO_SIGNED(602,11),
TO_SIGNED(629,11),
TO_SIGNED(653,11),
TO_SIGNED(675,11),
TO_SIGNED(694,11),
TO_SIGNED(711,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(729,11),
TO_SIGNED(716,11),
TO_SIGNED(701,11),
TO_SIGNED(683,11),
TO_SIGNED(662,11),
TO_SIGNED(639,11),
TO_SIGNED(613,11),
TO_SIGNED(584,11),
TO_SIGNED(554,11),
TO_SIGNED(521,11),
TO_SIGNED(486,11),
TO_SIGNED(449,11),
TO_SIGNED(411,11),
TO_SIGNED(371,11),
TO_SIGNED(329,11),
TO_SIGNED(286,11),
TO_SIGNED(242,11),
TO_SIGNED(197,11),
TO_SIGNED(152,11),
TO_SIGNED(105,11),
TO_SIGNED(59,11),
TO_SIGNED(12,11),
TO_SIGNED(-35,11),
TO_SIGNED(-82,11),
TO_SIGNED(-129,11),
TO_SIGNED(-175,11),
TO_SIGNED(-220,11),
TO_SIGNED(-265,11),
TO_SIGNED(-308,11),
TO_SIGNED(-350,11),
TO_SIGNED(-391,11),
TO_SIGNED(-430,11),
TO_SIGNED(-468,11),
TO_SIGNED(-504,11),
TO_SIGNED(-538,11),
TO_SIGNED(-569,11),
TO_SIGNED(-599,11),
TO_SIGNED(-626,11),
TO_SIGNED(-651,11),
TO_SIGNED(-673,11),
TO_SIGNED(-692,11),
TO_SIGNED(-709,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-685,11),
TO_SIGNED(-664,11),
TO_SIGNED(-641,11),
TO_SIGNED(-616,11),
TO_SIGNED(-588,11),
TO_SIGNED(-557,11),
TO_SIGNED(-525,11),
TO_SIGNED(-490,11),
TO_SIGNED(-454,11),
TO_SIGNED(-415,11),
TO_SIGNED(-375,11),
TO_SIGNED(-334,11),
TO_SIGNED(-291,11),
TO_SIGNED(-247,11),
TO_SIGNED(-203,11),
TO_SIGNED(-157,11),
TO_SIGNED(-111,11),
TO_SIGNED(-64,11),
TO_SIGNED(-17,11),
TO_SIGNED(30,11),
TO_SIGNED(77,11),
TO_SIGNED(123,11),
TO_SIGNED(169,11),
TO_SIGNED(215,11),
TO_SIGNED(260,11),
TO_SIGNED(303,11),
TO_SIGNED(345,11),
TO_SIGNED(387,11),
TO_SIGNED(426,11),
TO_SIGNED(464,11),
TO_SIGNED(500,11),
TO_SIGNED(534,11),
TO_SIGNED(566,11),
TO_SIGNED(596,11),
TO_SIGNED(623,11),
TO_SIGNED(648,11),
TO_SIGNED(670,11),
TO_SIGNED(690,11),
TO_SIGNED(707,11),
TO_SIGNED(721,11),
TO_SIGNED(733,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(705,11),
TO_SIGNED(687,11),
TO_SIGNED(667,11),
TO_SIGNED(644,11),
TO_SIGNED(619,11),
TO_SIGNED(591,11),
TO_SIGNED(561,11),
TO_SIGNED(529,11),
TO_SIGNED(494,11),
TO_SIGNED(458,11),
TO_SIGNED(420,11),
TO_SIGNED(380,11),
TO_SIGNED(339,11),
TO_SIGNED(296,11),
TO_SIGNED(252,11),
TO_SIGNED(208,11),
TO_SIGNED(162,11),
TO_SIGNED(116,11),
TO_SIGNED(69,11),
TO_SIGNED(22,11),
TO_SIGNED(-25,11),
TO_SIGNED(-71,11),
TO_SIGNED(-118,11),
TO_SIGNED(-164,11),
TO_SIGNED(-210,11),
TO_SIGNED(-255,11),
TO_SIGNED(-298,11),
TO_SIGNED(-341,11),
TO_SIGNED(-382,11),
TO_SIGNED(-422,11),
TO_SIGNED(-460,11),
TO_SIGNED(-496,11),
TO_SIGNED(-530,11),
TO_SIGNED(-562,11),
TO_SIGNED(-592,11),
TO_SIGNED(-620,11),
TO_SIGNED(-645,11),
TO_SIGNED(-668,11),
TO_SIGNED(-688,11),
TO_SIGNED(-705,11),
TO_SIGNED(-720,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-721,11),
TO_SIGNED(-706,11),
TO_SIGNED(-689,11),
TO_SIGNED(-669,11),
TO_SIGNED(-647,11),
TO_SIGNED(-622,11),
TO_SIGNED(-594,11),
TO_SIGNED(-564,11),
TO_SIGNED(-532,11),
TO_SIGNED(-498,11),
TO_SIGNED(-462,11),
TO_SIGNED(-424,11),
TO_SIGNED(-385,11),
TO_SIGNED(-344,11),
TO_SIGNED(-301,11),
TO_SIGNED(-258,11),
TO_SIGNED(-213,11),
TO_SIGNED(-167,11),
TO_SIGNED(-121,11),
TO_SIGNED(-75,11),
TO_SIGNED(-28,11),
TO_SIGNED(19,11),
TO_SIGNED(66,11),
TO_SIGNED(113,11),
TO_SIGNED(159,11),
TO_SIGNED(205,11),
TO_SIGNED(249,11),
TO_SIGNED(293,11),
TO_SIGNED(336,11),
TO_SIGNED(377,11),
TO_SIGNED(417,11),
TO_SIGNED(455,11),
TO_SIGNED(492,11),
TO_SIGNED(526,11),
TO_SIGNED(559,11),
TO_SIGNED(589,11),
TO_SIGNED(617,11),
TO_SIGNED(642,11),
TO_SIGNED(665,11),
TO_SIGNED(686,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(708,11),
TO_SIGNED(691,11),
TO_SIGNED(672,11),
TO_SIGNED(650,11),
TO_SIGNED(625,11),
TO_SIGNED(598,11),
TO_SIGNED(568,11),
TO_SIGNED(536,11),
TO_SIGNED(502,11),
TO_SIGNED(466,11),
TO_SIGNED(429,11),
TO_SIGNED(389,11),
TO_SIGNED(348,11),
TO_SIGNED(306,11),
TO_SIGNED(263,11),
TO_SIGNED(218,11),
TO_SIGNED(173,11),
TO_SIGNED(127,11),
TO_SIGNED(80,11),
TO_SIGNED(33,11),
TO_SIGNED(-14,11),
TO_SIGNED(-61,11),
TO_SIGNED(-108,11),
TO_SIGNED(-154,11),
TO_SIGNED(-200,11),
TO_SIGNED(-244,11),
TO_SIGNED(-288,11),
TO_SIGNED(-331,11),
TO_SIGNED(-373,11),
TO_SIGNED(-413,11),
TO_SIGNED(-451,11),
TO_SIGNED(-488,11),
TO_SIGNED(-523,11),
TO_SIGNED(-555,11),
TO_SIGNED(-586,11),
TO_SIGNED(-614,11),
TO_SIGNED(-640,11),
TO_SIGNED(-663,11),
TO_SIGNED(-684,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-729,11),
TO_SIGNED(-739,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-710,11),
TO_SIGNED(-693,11),
TO_SIGNED(-674,11),
TO_SIGNED(-652,11),
TO_SIGNED(-628,11),
TO_SIGNED(-601,11),
TO_SIGNED(-571,11),
TO_SIGNED(-540,11),
TO_SIGNED(-506,11),
TO_SIGNED(-471,11),
TO_SIGNED(-433,11),
TO_SIGNED(-394,11),
TO_SIGNED(-353,11),
TO_SIGNED(-311,11),
TO_SIGNED(-268,11),
TO_SIGNED(-223,11),
TO_SIGNED(-178,11),
TO_SIGNED(-132,11),
TO_SIGNED(-85,11),
TO_SIGNED(-38,11),
TO_SIGNED(9,11),
TO_SIGNED(56,11),
TO_SIGNED(102,11),
TO_SIGNED(149,11),
TO_SIGNED(194,11),
TO_SIGNED(239,11),
TO_SIGNED(283,11),
TO_SIGNED(326,11),
TO_SIGNED(368,11),
TO_SIGNED(408,11),
TO_SIGNED(447,11),
TO_SIGNED(484,11),
TO_SIGNED(519,11),
TO_SIGNED(552,11),
TO_SIGNED(582,11),
TO_SIGNED(611,11),
TO_SIGNED(637,11),
TO_SIGNED(660,11),
TO_SIGNED(681,11),
TO_SIGNED(700,11),
TO_SIGNED(715,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(736,11),
TO_SIGNED(725,11),
TO_SIGNED(712,11),
TO_SIGNED(695,11),
TO_SIGNED(676,11),
TO_SIGNED(655,11),
TO_SIGNED(631,11),
TO_SIGNED(604,11),
TO_SIGNED(575,11),
TO_SIGNED(544,11),
TO_SIGNED(510,11),
TO_SIGNED(475,11),
TO_SIGNED(437,11),
TO_SIGNED(398,11),
TO_SIGNED(358,11),
TO_SIGNED(316,11),
TO_SIGNED(273,11),
TO_SIGNED(228,11),
TO_SIGNED(183,11),
TO_SIGNED(137,11),
TO_SIGNED(91,11),
TO_SIGNED(44,11),
TO_SIGNED(-3,11),
TO_SIGNED(-50,11),
TO_SIGNED(-97,11),
TO_SIGNED(-143,11),
TO_SIGNED(-189,11),
TO_SIGNED(-234,11),
TO_SIGNED(-278,11),
TO_SIGNED(-322,11),
TO_SIGNED(-363,11),
TO_SIGNED(-404,11),
TO_SIGNED(-443,11),
TO_SIGNED(-480,11),
TO_SIGNED(-515,11),
TO_SIGNED(-548,11),
TO_SIGNED(-579,11),
TO_SIGNED(-608,11),
TO_SIGNED(-634,11),
TO_SIGNED(-658,11),
TO_SIGNED(-679,11),
TO_SIGNED(-698,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-679,11),
TO_SIGNED(-657,11),
TO_SIGNED(-633,11),
TO_SIGNED(-607,11),
TO_SIGNED(-578,11),
TO_SIGNED(-547,11),
TO_SIGNED(-514,11),
TO_SIGNED(-479,11),
TO_SIGNED(-442,11),
TO_SIGNED(-403,11),
TO_SIGNED(-362,11),
TO_SIGNED(-321,11),
TO_SIGNED(-277,11),
TO_SIGNED(-233,11),
TO_SIGNED(-188,11),
TO_SIGNED(-142,11),
TO_SIGNED(-96,11),
TO_SIGNED(-49,11),
TO_SIGNED(-2,11),
TO_SIGNED(45,11),
TO_SIGNED(92,11),
TO_SIGNED(138,11),
TO_SIGNED(184,11),
TO_SIGNED(229,11),
TO_SIGNED(274,11),
TO_SIGNED(317,11),
TO_SIGNED(359,11),
TO_SIGNED(399,11),
TO_SIGNED(438,11),
TO_SIGNED(476,11),
TO_SIGNED(511,11),
TO_SIGNED(544,11),
TO_SIGNED(576,11),
TO_SIGNED(605,11),
TO_SIGNED(631,11),
TO_SIGNED(655,11),
TO_SIGNED(677,11),
TO_SIGNED(696,11),
TO_SIGNED(712,11),
TO_SIGNED(725,11),
TO_SIGNED(736,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(715,11),
TO_SIGNED(699,11),
TO_SIGNED(681,11),
TO_SIGNED(660,11),
TO_SIGNED(636,11),
TO_SIGNED(610,11),
TO_SIGNED(582,11),
TO_SIGNED(551,11),
TO_SIGNED(518,11),
TO_SIGNED(483,11),
TO_SIGNED(446,11),
TO_SIGNED(407,11),
TO_SIGNED(367,11),
TO_SIGNED(325,11),
TO_SIGNED(282,11),
TO_SIGNED(238,11),
TO_SIGNED(193,11),
TO_SIGNED(148,11),
TO_SIGNED(101,11),
TO_SIGNED(54,11),
TO_SIGNED(7,11),
TO_SIGNED(-40,11),
TO_SIGNED(-86,11),
TO_SIGNED(-133,11),
TO_SIGNED(-179,11),
TO_SIGNED(-224,11),
TO_SIGNED(-269,11),
TO_SIGNED(-312,11),
TO_SIGNED(-354,11),
TO_SIGNED(-395,11),
TO_SIGNED(-434,11),
TO_SIGNED(-471,11),
TO_SIGNED(-507,11),
TO_SIGNED(-541,11),
TO_SIGNED(-572,11),
TO_SIGNED(-601,11),
TO_SIGNED(-628,11),
TO_SIGNED(-653,11),
TO_SIGNED(-675,11),
TO_SIGNED(-694,11),
TO_SIGNED(-710,11),
TO_SIGNED(-724,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-701,11),
TO_SIGNED(-683,11),
TO_SIGNED(-662,11),
TO_SIGNED(-639,11),
TO_SIGNED(-613,11),
TO_SIGNED(-585,11),
TO_SIGNED(-554,11),
TO_SIGNED(-522,11),
TO_SIGNED(-487,11),
TO_SIGNED(-450,11),
TO_SIGNED(-412,11),
TO_SIGNED(-372,11),
TO_SIGNED(-330,11),
TO_SIGNED(-287,11),
TO_SIGNED(-243,11),
TO_SIGNED(-198,11),
TO_SIGNED(-153,11),
TO_SIGNED(-106,11),
TO_SIGNED(-60,11),
TO_SIGNED(-13,11),
TO_SIGNED(34,11),
TO_SIGNED(81,11),
TO_SIGNED(128,11),
TO_SIGNED(174,11),
TO_SIGNED(219,11),
TO_SIGNED(264,11),
TO_SIGNED(307,11),
TO_SIGNED(349,11),
TO_SIGNED(390,11),
TO_SIGNED(430,11),
TO_SIGNED(467,11),
TO_SIGNED(503,11),
TO_SIGNED(537,11),
TO_SIGNED(569,11),
TO_SIGNED(598,11),
TO_SIGNED(625,11),
TO_SIGNED(650,11),
TO_SIGNED(672,11),
TO_SIGNED(692,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(730,11),
TO_SIGNED(718,11),
TO_SIGNED(703,11),
TO_SIGNED(685,11),
TO_SIGNED(665,11),
TO_SIGNED(642,11),
TO_SIGNED(616,11),
TO_SIGNED(588,11),
TO_SIGNED(558,11),
TO_SIGNED(526,11),
TO_SIGNED(491,11),
TO_SIGNED(455,11),
TO_SIGNED(416,11),
TO_SIGNED(376,11),
TO_SIGNED(335,11),
TO_SIGNED(292,11),
TO_SIGNED(248,11),
TO_SIGNED(204,11),
TO_SIGNED(158,11),
TO_SIGNED(112,11),
TO_SIGNED(65,11),
TO_SIGNED(18,11),
TO_SIGNED(-29,11),
TO_SIGNED(-76,11),
TO_SIGNED(-122,11),
TO_SIGNED(-168,11),
TO_SIGNED(-214,11),
TO_SIGNED(-259,11),
TO_SIGNED(-302,11),
TO_SIGNED(-345,11),
TO_SIGNED(-386,11),
TO_SIGNED(-425,11),
TO_SIGNED(-463,11),
TO_SIGNED(-499,11),
TO_SIGNED(-533,11),
TO_SIGNED(-565,11),
TO_SIGNED(-595,11),
TO_SIGNED(-622,11),
TO_SIGNED(-647,11),
TO_SIGNED(-670,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-721,11),
TO_SIGNED(-733,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-720,11),
TO_SIGNED(-705,11),
TO_SIGNED(-688,11),
TO_SIGNED(-667,11),
TO_SIGNED(-645,11),
TO_SIGNED(-619,11),
TO_SIGNED(-592,11),
TO_SIGNED(-562,11),
TO_SIGNED(-529,11),
TO_SIGNED(-495,11),
TO_SIGNED(-459,11),
TO_SIGNED(-421,11),
TO_SIGNED(-381,11),
TO_SIGNED(-340,11),
TO_SIGNED(-297,11),
TO_SIGNED(-254,11),
TO_SIGNED(-209,11),
TO_SIGNED(-163,11),
TO_SIGNED(-117,11),
TO_SIGNED(-70,11),
TO_SIGNED(-24,11),
TO_SIGNED(24,11),
TO_SIGNED(70,11),
TO_SIGNED(117,11),
TO_SIGNED(163,11),
TO_SIGNED(209,11),
TO_SIGNED(254,11),
TO_SIGNED(297,11),
TO_SIGNED(340,11),
TO_SIGNED(381,11),
TO_SIGNED(421,11),
TO_SIGNED(459,11),
TO_SIGNED(495,11),
TO_SIGNED(529,11),
TO_SIGNED(562,11),
TO_SIGNED(592,11),
TO_SIGNED(619,11),
TO_SIGNED(645,11),
TO_SIGNED(667,11),
TO_SIGNED(688,11),
TO_SIGNED(705,11),
TO_SIGNED(720,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(733,11),
TO_SIGNED(721,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(670,11),
TO_SIGNED(647,11),
TO_SIGNED(622,11),
TO_SIGNED(595,11),
TO_SIGNED(565,11),
TO_SIGNED(533,11),
TO_SIGNED(499,11),
TO_SIGNED(463,11),
TO_SIGNED(425,11),
TO_SIGNED(386,11),
TO_SIGNED(345,11),
TO_SIGNED(302,11),
TO_SIGNED(259,11),
TO_SIGNED(214,11),
TO_SIGNED(168,11),
TO_SIGNED(122,11),
TO_SIGNED(76,11),
TO_SIGNED(29,11),
TO_SIGNED(-18,11),
TO_SIGNED(-65,11),
TO_SIGNED(-112,11),
TO_SIGNED(-158,11),
TO_SIGNED(-204,11),
TO_SIGNED(-248,11),
TO_SIGNED(-292,11),
TO_SIGNED(-335,11),
TO_SIGNED(-376,11),
TO_SIGNED(-416,11),
TO_SIGNED(-455,11),
TO_SIGNED(-491,11),
TO_SIGNED(-526,11),
TO_SIGNED(-558,11),
TO_SIGNED(-588,11),
TO_SIGNED(-616,11),
TO_SIGNED(-642,11),
TO_SIGNED(-665,11),
TO_SIGNED(-685,11),
TO_SIGNED(-703,11),
TO_SIGNED(-718,11),
TO_SIGNED(-730,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-692,11),
TO_SIGNED(-672,11),
TO_SIGNED(-650,11),
TO_SIGNED(-625,11),
TO_SIGNED(-598,11),
TO_SIGNED(-569,11),
TO_SIGNED(-537,11),
TO_SIGNED(-503,11),
TO_SIGNED(-467,11),
TO_SIGNED(-430,11),
TO_SIGNED(-390,11),
TO_SIGNED(-349,11),
TO_SIGNED(-307,11),
TO_SIGNED(-264,11),
TO_SIGNED(-219,11),
TO_SIGNED(-174,11),
TO_SIGNED(-128,11),
TO_SIGNED(-81,11),
TO_SIGNED(-34,11),
TO_SIGNED(13,11),
TO_SIGNED(60,11),
TO_SIGNED(106,11),
TO_SIGNED(153,11),
TO_SIGNED(198,11),
TO_SIGNED(243,11),
TO_SIGNED(287,11),
TO_SIGNED(330,11),
TO_SIGNED(372,11),
TO_SIGNED(412,11),
TO_SIGNED(450,11),
TO_SIGNED(487,11),
TO_SIGNED(522,11),
TO_SIGNED(554,11),
TO_SIGNED(585,11),
TO_SIGNED(613,11),
TO_SIGNED(639,11),
TO_SIGNED(662,11),
TO_SIGNED(683,11),
TO_SIGNED(701,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(724,11),
TO_SIGNED(710,11),
TO_SIGNED(694,11),
TO_SIGNED(675,11),
TO_SIGNED(653,11),
TO_SIGNED(628,11),
TO_SIGNED(601,11),
TO_SIGNED(572,11),
TO_SIGNED(541,11),
TO_SIGNED(507,11),
TO_SIGNED(471,11),
TO_SIGNED(434,11),
TO_SIGNED(395,11),
TO_SIGNED(354,11),
TO_SIGNED(312,11),
TO_SIGNED(269,11),
TO_SIGNED(224,11),
TO_SIGNED(179,11),
TO_SIGNED(133,11),
TO_SIGNED(86,11),
TO_SIGNED(40,11),
TO_SIGNED(-7,11),
TO_SIGNED(-54,11),
TO_SIGNED(-101,11),
TO_SIGNED(-148,11),
TO_SIGNED(-193,11),
TO_SIGNED(-238,11),
TO_SIGNED(-282,11),
TO_SIGNED(-325,11),
TO_SIGNED(-367,11),
TO_SIGNED(-407,11),
TO_SIGNED(-446,11),
TO_SIGNED(-483,11),
TO_SIGNED(-518,11),
TO_SIGNED(-551,11),
TO_SIGNED(-582,11),
TO_SIGNED(-610,11),
TO_SIGNED(-636,11),
TO_SIGNED(-660,11),
TO_SIGNED(-681,11),
TO_SIGNED(-699,11),
TO_SIGNED(-715,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-736,11),
TO_SIGNED(-725,11),
TO_SIGNED(-712,11),
TO_SIGNED(-696,11),
TO_SIGNED(-677,11),
TO_SIGNED(-655,11),
TO_SIGNED(-631,11),
TO_SIGNED(-605,11),
TO_SIGNED(-576,11),
TO_SIGNED(-544,11),
TO_SIGNED(-511,11),
TO_SIGNED(-476,11),
TO_SIGNED(-438,11),
TO_SIGNED(-399,11),
TO_SIGNED(-359,11),
TO_SIGNED(-317,11),
TO_SIGNED(-274,11),
TO_SIGNED(-229,11),
TO_SIGNED(-184,11),
TO_SIGNED(-138,11),
TO_SIGNED(-92,11),
TO_SIGNED(-45,11),
TO_SIGNED(2,11),
TO_SIGNED(49,11),
TO_SIGNED(96,11),
TO_SIGNED(142,11),
TO_SIGNED(188,11),
TO_SIGNED(233,11),
TO_SIGNED(277,11),
TO_SIGNED(321,11),
TO_SIGNED(362,11),
TO_SIGNED(403,11),
TO_SIGNED(442,11),
TO_SIGNED(479,11),
TO_SIGNED(514,11),
TO_SIGNED(547,11),
TO_SIGNED(578,11),
TO_SIGNED(607,11),
TO_SIGNED(633,11),
TO_SIGNED(657,11),
TO_SIGNED(679,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(698,11),
TO_SIGNED(679,11),
TO_SIGNED(658,11),
TO_SIGNED(634,11),
TO_SIGNED(608,11),
TO_SIGNED(579,11),
TO_SIGNED(548,11),
TO_SIGNED(515,11),
TO_SIGNED(480,11),
TO_SIGNED(443,11),
TO_SIGNED(404,11),
TO_SIGNED(363,11),
TO_SIGNED(322,11),
TO_SIGNED(278,11),
TO_SIGNED(234,11),
TO_SIGNED(189,11),
TO_SIGNED(143,11),
TO_SIGNED(97,11),
TO_SIGNED(50,11),
TO_SIGNED(3,11),
TO_SIGNED(-44,11),
TO_SIGNED(-91,11),
TO_SIGNED(-137,11),
TO_SIGNED(-183,11),
TO_SIGNED(-228,11),
TO_SIGNED(-273,11),
TO_SIGNED(-316,11),
TO_SIGNED(-358,11),
TO_SIGNED(-398,11),
TO_SIGNED(-437,11),
TO_SIGNED(-475,11),
TO_SIGNED(-510,11),
TO_SIGNED(-544,11),
TO_SIGNED(-575,11),
TO_SIGNED(-604,11),
TO_SIGNED(-631,11),
TO_SIGNED(-655,11),
TO_SIGNED(-676,11),
TO_SIGNED(-695,11),
TO_SIGNED(-712,11),
TO_SIGNED(-725,11),
TO_SIGNED(-736,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-715,11),
TO_SIGNED(-700,11),
TO_SIGNED(-681,11),
TO_SIGNED(-660,11),
TO_SIGNED(-637,11),
TO_SIGNED(-611,11),
TO_SIGNED(-582,11),
TO_SIGNED(-552,11),
TO_SIGNED(-519,11),
TO_SIGNED(-484,11),
TO_SIGNED(-447,11),
TO_SIGNED(-408,11),
TO_SIGNED(-368,11),
TO_SIGNED(-326,11),
TO_SIGNED(-283,11),
TO_SIGNED(-239,11),
TO_SIGNED(-194,11),
TO_SIGNED(-149,11),
TO_SIGNED(-102,11),
TO_SIGNED(-56,11),
TO_SIGNED(-9,11),
TO_SIGNED(38,11),
TO_SIGNED(85,11),
TO_SIGNED(132,11),
TO_SIGNED(178,11),
TO_SIGNED(223,11),
TO_SIGNED(268,11),
TO_SIGNED(311,11),
TO_SIGNED(353,11),
TO_SIGNED(394,11),
TO_SIGNED(433,11),
TO_SIGNED(471,11),
TO_SIGNED(506,11),
TO_SIGNED(540,11),
TO_SIGNED(571,11),
TO_SIGNED(601,11),
TO_SIGNED(628,11),
TO_SIGNED(652,11),
TO_SIGNED(674,11),
TO_SIGNED(693,11),
TO_SIGNED(710,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(739,11),
TO_SIGNED(729,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(684,11),
TO_SIGNED(663,11),
TO_SIGNED(640,11),
TO_SIGNED(614,11),
TO_SIGNED(586,11),
TO_SIGNED(555,11),
TO_SIGNED(523,11),
TO_SIGNED(488,11),
TO_SIGNED(451,11),
TO_SIGNED(413,11),
TO_SIGNED(373,11),
TO_SIGNED(331,11),
TO_SIGNED(288,11),
TO_SIGNED(244,11),
TO_SIGNED(200,11),
TO_SIGNED(154,11),
TO_SIGNED(108,11),
TO_SIGNED(61,11),
TO_SIGNED(14,11),
TO_SIGNED(-33,11),
TO_SIGNED(-80,11),
TO_SIGNED(-127,11),
TO_SIGNED(-173,11),
TO_SIGNED(-218,11),
TO_SIGNED(-263,11),
TO_SIGNED(-306,11),
TO_SIGNED(-348,11),
TO_SIGNED(-389,11),
TO_SIGNED(-429,11),
TO_SIGNED(-466,11),
TO_SIGNED(-502,11),
TO_SIGNED(-536,11),
TO_SIGNED(-568,11),
TO_SIGNED(-598,11),
TO_SIGNED(-625,11),
TO_SIGNED(-650,11),
TO_SIGNED(-672,11),
TO_SIGNED(-691,11),
TO_SIGNED(-708,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-686,11),
TO_SIGNED(-665,11),
TO_SIGNED(-642,11),
TO_SIGNED(-617,11),
TO_SIGNED(-589,11),
TO_SIGNED(-559,11),
TO_SIGNED(-526,11),
TO_SIGNED(-492,11),
TO_SIGNED(-455,11),
TO_SIGNED(-417,11),
TO_SIGNED(-377,11),
TO_SIGNED(-336,11),
TO_SIGNED(-293,11),
TO_SIGNED(-249,11),
TO_SIGNED(-205,11),
TO_SIGNED(-159,11),
TO_SIGNED(-113,11),
TO_SIGNED(-66,11),
TO_SIGNED(-19,11),
TO_SIGNED(28,11),
TO_SIGNED(75,11),
TO_SIGNED(121,11),
TO_SIGNED(167,11),
TO_SIGNED(213,11),
TO_SIGNED(258,11),
TO_SIGNED(301,11),
TO_SIGNED(344,11),
TO_SIGNED(385,11),
TO_SIGNED(424,11),
TO_SIGNED(462,11),
TO_SIGNED(498,11),
TO_SIGNED(532,11),
TO_SIGNED(564,11),
TO_SIGNED(594,11),
TO_SIGNED(622,11),
TO_SIGNED(647,11),
TO_SIGNED(669,11),
TO_SIGNED(689,11),
TO_SIGNED(706,11),
TO_SIGNED(721,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(720,11),
TO_SIGNED(705,11),
TO_SIGNED(688,11),
TO_SIGNED(668,11),
TO_SIGNED(645,11),
TO_SIGNED(620,11),
TO_SIGNED(592,11),
TO_SIGNED(562,11),
TO_SIGNED(530,11),
TO_SIGNED(496,11),
TO_SIGNED(460,11),
TO_SIGNED(422,11),
TO_SIGNED(382,11),
TO_SIGNED(341,11),
TO_SIGNED(298,11),
TO_SIGNED(255,11),
TO_SIGNED(210,11),
TO_SIGNED(164,11),
TO_SIGNED(118,11),
TO_SIGNED(71,11),
TO_SIGNED(25,11),
TO_SIGNED(-22,11),
TO_SIGNED(-69,11),
TO_SIGNED(-116,11),
TO_SIGNED(-162,11),
TO_SIGNED(-208,11),
TO_SIGNED(-252,11),
TO_SIGNED(-296,11),
TO_SIGNED(-339,11),
TO_SIGNED(-380,11),
TO_SIGNED(-420,11),
TO_SIGNED(-458,11),
TO_SIGNED(-494,11),
TO_SIGNED(-529,11),
TO_SIGNED(-561,11),
TO_SIGNED(-591,11),
TO_SIGNED(-619,11),
TO_SIGNED(-644,11),
TO_SIGNED(-667,11),
TO_SIGNED(-687,11),
TO_SIGNED(-705,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-733,11),
TO_SIGNED(-721,11),
TO_SIGNED(-707,11),
TO_SIGNED(-690,11),
TO_SIGNED(-670,11),
TO_SIGNED(-648,11),
TO_SIGNED(-623,11),
TO_SIGNED(-596,11),
TO_SIGNED(-566,11),
TO_SIGNED(-534,11),
TO_SIGNED(-500,11),
TO_SIGNED(-464,11),
TO_SIGNED(-426,11),
TO_SIGNED(-387,11),
TO_SIGNED(-345,11),
TO_SIGNED(-303,11),
TO_SIGNED(-260,11),
TO_SIGNED(-215,11),
TO_SIGNED(-169,11),
TO_SIGNED(-123,11),
TO_SIGNED(-77,11),
TO_SIGNED(-30,11),
TO_SIGNED(17,11),
TO_SIGNED(64,11),
TO_SIGNED(111,11),
TO_SIGNED(157,11),
TO_SIGNED(203,11),
TO_SIGNED(247,11),
TO_SIGNED(291,11),
TO_SIGNED(334,11),
TO_SIGNED(375,11),
TO_SIGNED(415,11),
TO_SIGNED(454,11),
TO_SIGNED(490,11),
TO_SIGNED(525,11),
TO_SIGNED(557,11),
TO_SIGNED(588,11),
TO_SIGNED(616,11),
TO_SIGNED(641,11),
TO_SIGNED(664,11),
TO_SIGNED(685,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(709,11),
TO_SIGNED(692,11),
TO_SIGNED(673,11),
TO_SIGNED(651,11),
TO_SIGNED(626,11),
TO_SIGNED(599,11),
TO_SIGNED(569,11),
TO_SIGNED(538,11),
TO_SIGNED(504,11),
TO_SIGNED(468,11),
TO_SIGNED(430,11),
TO_SIGNED(391,11),
TO_SIGNED(350,11),
TO_SIGNED(308,11),
TO_SIGNED(265,11),
TO_SIGNED(220,11),
TO_SIGNED(175,11),
TO_SIGNED(129,11),
TO_SIGNED(82,11),
TO_SIGNED(35,11),
TO_SIGNED(-12,11),
TO_SIGNED(-59,11),
TO_SIGNED(-105,11),
TO_SIGNED(-152,11),
TO_SIGNED(-197,11),
TO_SIGNED(-242,11),
TO_SIGNED(-286,11),
TO_SIGNED(-329,11),
TO_SIGNED(-371,11),
TO_SIGNED(-411,11),
TO_SIGNED(-449,11),
TO_SIGNED(-486,11),
TO_SIGNED(-521,11),
TO_SIGNED(-554,11),
TO_SIGNED(-584,11),
TO_SIGNED(-613,11),
TO_SIGNED(-639,11),
TO_SIGNED(-662,11),
TO_SIGNED(-683,11),
TO_SIGNED(-701,11),
TO_SIGNED(-716,11),
TO_SIGNED(-729,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-711,11),
TO_SIGNED(-694,11),
TO_SIGNED(-675,11),
TO_SIGNED(-653,11),
TO_SIGNED(-629,11),
TO_SIGNED(-602,11),
TO_SIGNED(-573,11),
TO_SIGNED(-541,11),
TO_SIGNED(-508,11),
TO_SIGNED(-472,11),
TO_SIGNED(-435,11),
TO_SIGNED(-396,11),
TO_SIGNED(-355,11),
TO_SIGNED(-313,11),
TO_SIGNED(-270,11),
TO_SIGNED(-225,11),
TO_SIGNED(-180,11),
TO_SIGNED(-134,11),
TO_SIGNED(-87,11),
TO_SIGNED(-41,11),
TO_SIGNED(6,11),
TO_SIGNED(53,11),
TO_SIGNED(100,11),
TO_SIGNED(147,11),
TO_SIGNED(192,11),
TO_SIGNED(237,11),
TO_SIGNED(281,11),
TO_SIGNED(324,11),
TO_SIGNED(366,11),
TO_SIGNED(406,11),
TO_SIGNED(445,11),
TO_SIGNED(482,11),
TO_SIGNED(517,11),
TO_SIGNED(550,11),
TO_SIGNED(581,11),
TO_SIGNED(610,11),
TO_SIGNED(636,11),
TO_SIGNED(659,11),
TO_SIGNED(681,11),
TO_SIGNED(699,11),
TO_SIGNED(715,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(712,11),
TO_SIGNED(696,11),
TO_SIGNED(677,11),
TO_SIGNED(656,11),
TO_SIGNED(632,11),
TO_SIGNED(605,11),
TO_SIGNED(576,11),
TO_SIGNED(545,11),
TO_SIGNED(512,11),
TO_SIGNED(476,11),
TO_SIGNED(439,11),
TO_SIGNED(400,11),
TO_SIGNED(360,11),
TO_SIGNED(318,11),
TO_SIGNED(275,11),
TO_SIGNED(230,11),
TO_SIGNED(185,11),
TO_SIGNED(139,11),
TO_SIGNED(93,11),
TO_SIGNED(46,11),
TO_SIGNED(-1,11),
TO_SIGNED(-48,11),
TO_SIGNED(-95,11),
TO_SIGNED(-141,11),
TO_SIGNED(-187,11),
TO_SIGNED(-232,11),
TO_SIGNED(-276,11),
TO_SIGNED(-320,11),
TO_SIGNED(-362,11),
TO_SIGNED(-402,11),
TO_SIGNED(-441,11),
TO_SIGNED(-478,11),
TO_SIGNED(-513,11),
TO_SIGNED(-547,11),
TO_SIGNED(-578,11),
TO_SIGNED(-606,11),
TO_SIGNED(-633,11),
TO_SIGNED(-657,11),
TO_SIGNED(-678,11),
TO_SIGNED(-697,11),
TO_SIGNED(-713,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-714,11),
TO_SIGNED(-698,11),
TO_SIGNED(-680,11),
TO_SIGNED(-658,11),
TO_SIGNED(-635,11),
TO_SIGNED(-608,11),
TO_SIGNED(-580,11),
TO_SIGNED(-549,11),
TO_SIGNED(-516,11),
TO_SIGNED(-480,11),
TO_SIGNED(-443,11),
TO_SIGNED(-405,11),
TO_SIGNED(-364,11),
TO_SIGNED(-323,11),
TO_SIGNED(-279,11),
TO_SIGNED(-235,11),
TO_SIGNED(-190,11),
TO_SIGNED(-144,11),
TO_SIGNED(-98,11),
TO_SIGNED(-51,11),
TO_SIGNED(-4,11),
TO_SIGNED(43,11),
TO_SIGNED(90,11),
TO_SIGNED(136,11),
TO_SIGNED(182,11),
TO_SIGNED(227,11),
TO_SIGNED(272,11),
TO_SIGNED(315,11),
TO_SIGNED(357,11),
TO_SIGNED(397,11),
TO_SIGNED(437,11),
TO_SIGNED(474,11),
TO_SIGNED(509,11),
TO_SIGNED(543,11),
TO_SIGNED(574,11),
TO_SIGNED(603,11),
TO_SIGNED(630,11),
TO_SIGNED(654,11),
TO_SIGNED(676,11),
TO_SIGNED(695,11),
TO_SIGNED(711,11),
TO_SIGNED(725,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(716,11),
TO_SIGNED(700,11),
TO_SIGNED(682,11),
TO_SIGNED(661,11),
TO_SIGNED(637,11),
TO_SIGNED(611,11),
TO_SIGNED(583,11),
TO_SIGNED(552,11),
TO_SIGNED(519,11),
TO_SIGNED(485,11),
TO_SIGNED(448,11),
TO_SIGNED(409,11),
TO_SIGNED(369,11),
TO_SIGNED(327,11),
TO_SIGNED(284,11),
TO_SIGNED(240,11),
TO_SIGNED(195,11),
TO_SIGNED(150,11),
TO_SIGNED(103,11),
TO_SIGNED(57,11),
TO_SIGNED(10,11),
TO_SIGNED(-37,11),
TO_SIGNED(-84,11),
TO_SIGNED(-131,11),
TO_SIGNED(-177,11),
TO_SIGNED(-222,11),
TO_SIGNED(-267,11),
TO_SIGNED(-310,11),
TO_SIGNED(-352,11),
TO_SIGNED(-393,11),
TO_SIGNED(-432,11),
TO_SIGNED(-470,11),
TO_SIGNED(-505,11),
TO_SIGNED(-539,11),
TO_SIGNED(-571,11),
TO_SIGNED(-600,11),
TO_SIGNED(-627,11),
TO_SIGNED(-652,11),
TO_SIGNED(-674,11),
TO_SIGNED(-693,11),
TO_SIGNED(-710,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-702,11),
TO_SIGNED(-684,11),
TO_SIGNED(-663,11),
TO_SIGNED(-640,11),
TO_SIGNED(-615,11),
TO_SIGNED(-586,11),
TO_SIGNED(-556,11),
TO_SIGNED(-523,11),
TO_SIGNED(-489,11),
TO_SIGNED(-452,11),
TO_SIGNED(-414,11),
TO_SIGNED(-374,11),
TO_SIGNED(-332,11),
TO_SIGNED(-289,11),
TO_SIGNED(-245,11),
TO_SIGNED(-201,11),
TO_SIGNED(-155,11),
TO_SIGNED(-109,11),
TO_SIGNED(-62,11),
TO_SIGNED(-15,11),
TO_SIGNED(32,11),
TO_SIGNED(79,11),
TO_SIGNED(125,11),
TO_SIGNED(172,11),
TO_SIGNED(217,11),
TO_SIGNED(262,11),
TO_SIGNED(305,11),
TO_SIGNED(347,11),
TO_SIGNED(388,11),
TO_SIGNED(428,11),
TO_SIGNED(466,11),
TO_SIGNED(501,11),
TO_SIGNED(535,11),
TO_SIGNED(567,11),
TO_SIGNED(597,11),
TO_SIGNED(624,11),
TO_SIGNED(649,11),
TO_SIGNED(671,11),
TO_SIGNED(691,11),
TO_SIGNED(708,11),
TO_SIGNED(722,11),
TO_SIGNED(733,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(704,11),
TO_SIGNED(686,11),
TO_SIGNED(666,11),
TO_SIGNED(643,11),
TO_SIGNED(618,11),
TO_SIGNED(590,11),
TO_SIGNED(559,11),
TO_SIGNED(527,11),
TO_SIGNED(493,11),
TO_SIGNED(456,11),
TO_SIGNED(418,11),
TO_SIGNED(378,11),
TO_SIGNED(337,11),
TO_SIGNED(294,11),
TO_SIGNED(250,11),
TO_SIGNED(206,11),
TO_SIGNED(160,11),
TO_SIGNED(114,11),
TO_SIGNED(67,11),
TO_SIGNED(20,11),
TO_SIGNED(-27,11),
TO_SIGNED(-74,11),
TO_SIGNED(-120,11),
TO_SIGNED(-166,11),
TO_SIGNED(-212,11),
TO_SIGNED(-257,11),
TO_SIGNED(-300,11),
TO_SIGNED(-343,11),
TO_SIGNED(-384,11),
TO_SIGNED(-423,11),
TO_SIGNED(-461,11),
TO_SIGNED(-497,11),
TO_SIGNED(-532,11),
TO_SIGNED(-564,11),
TO_SIGNED(-594,11),
TO_SIGNED(-621,11),
TO_SIGNED(-646,11),
TO_SIGNED(-669,11),
TO_SIGNED(-689,11),
TO_SIGNED(-706,11),
TO_SIGNED(-721,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-720,11),
TO_SIGNED(-706,11),
TO_SIGNED(-688,11),
TO_SIGNED(-668,11),
TO_SIGNED(-646,11),
TO_SIGNED(-621,11),
TO_SIGNED(-593,11),
TO_SIGNED(-563,11),
TO_SIGNED(-531,11),
TO_SIGNED(-497,11),
TO_SIGNED(-460,11),
TO_SIGNED(-422,11),
TO_SIGNED(-383,11),
TO_SIGNED(-342,11),
TO_SIGNED(-299,11),
TO_SIGNED(-256,11),
TO_SIGNED(-211,11),
TO_SIGNED(-165,11),
TO_SIGNED(-119,11),
TO_SIGNED(-73,11),
TO_SIGNED(-26,11),
TO_SIGNED(21,11),
TO_SIGNED(68,11),
TO_SIGNED(115,11),
TO_SIGNED(161,11),
TO_SIGNED(207,11),
TO_SIGNED(251,11),
TO_SIGNED(295,11),
TO_SIGNED(338,11),
TO_SIGNED(379,11),
TO_SIGNED(419,11),
TO_SIGNED(457,11),
TO_SIGNED(493,11),
TO_SIGNED(528,11),
TO_SIGNED(560,11),
TO_SIGNED(590,11),
TO_SIGNED(618,11),
TO_SIGNED(644,11),
TO_SIGNED(666,11),
TO_SIGNED(687,11),
TO_SIGNED(704,11),
TO_SIGNED(719,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(671,11),
TO_SIGNED(648,11),
TO_SIGNED(624,11),
TO_SIGNED(596,11),
TO_SIGNED(567,11),
TO_SIGNED(535,11),
TO_SIGNED(501,11),
TO_SIGNED(465,11),
TO_SIGNED(427,11),
TO_SIGNED(387,11),
TO_SIGNED(346,11),
TO_SIGNED(304,11),
TO_SIGNED(261,11),
TO_SIGNED(216,11),
TO_SIGNED(171,11),
TO_SIGNED(124,11),
TO_SIGNED(78,11),
TO_SIGNED(31,11),
TO_SIGNED(-16,11),
TO_SIGNED(-63,11),
TO_SIGNED(-110,11),
TO_SIGNED(-156,11),
TO_SIGNED(-202,11),
TO_SIGNED(-246,11),
TO_SIGNED(-290,11),
TO_SIGNED(-333,11),
TO_SIGNED(-375,11),
TO_SIGNED(-415,11),
TO_SIGNED(-453,11),
TO_SIGNED(-489,11),
TO_SIGNED(-524,11),
TO_SIGNED(-557,11),
TO_SIGNED(-587,11),
TO_SIGNED(-615,11),
TO_SIGNED(-641,11),
TO_SIGNED(-664,11),
TO_SIGNED(-685,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-730,11),
TO_SIGNED(-739,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-693,11),
TO_SIGNED(-673,11),
TO_SIGNED(-651,11),
TO_SIGNED(-627,11),
TO_SIGNED(-599,11),
TO_SIGNED(-570,11),
TO_SIGNED(-538,11),
TO_SIGNED(-505,11),
TO_SIGNED(-469,11),
TO_SIGNED(-431,11),
TO_SIGNED(-392,11),
TO_SIGNED(-351,11),
TO_SIGNED(-309,11),
TO_SIGNED(-266,11),
TO_SIGNED(-221,11),
TO_SIGNED(-176,11),
TO_SIGNED(-130,11),
TO_SIGNED(-83,11),
TO_SIGNED(-36,11),
TO_SIGNED(11,11),
TO_SIGNED(58,11),
TO_SIGNED(104,11),
TO_SIGNED(151,11),
TO_SIGNED(196,11),
TO_SIGNED(241,11),
TO_SIGNED(285,11),
TO_SIGNED(328,11),
TO_SIGNED(370,11),
TO_SIGNED(410,11),
TO_SIGNED(449,11),
TO_SIGNED(485,11),
TO_SIGNED(520,11),
TO_SIGNED(553,11),
TO_SIGNED(584,11),
TO_SIGNED(612,11),
TO_SIGNED(638,11),
TO_SIGNED(661,11),
TO_SIGNED(682,11),
TO_SIGNED(700,11),
TO_SIGNED(716,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(725,11),
TO_SIGNED(711,11),
TO_SIGNED(695,11),
TO_SIGNED(675,11),
TO_SIGNED(654,11),
TO_SIGNED(629,11),
TO_SIGNED(603,11),
TO_SIGNED(574,11),
TO_SIGNED(542,11),
TO_SIGNED(509,11),
TO_SIGNED(473,11),
TO_SIGNED(436,11),
TO_SIGNED(397,11),
TO_SIGNED(356,11),
TO_SIGNED(314,11),
TO_SIGNED(271,11),
TO_SIGNED(226,11),
TO_SIGNED(181,11),
TO_SIGNED(135,11),
TO_SIGNED(88,11),
TO_SIGNED(42,11),
TO_SIGNED(-5,11),
TO_SIGNED(-52,11),
TO_SIGNED(-99,11),
TO_SIGNED(-145,11),
TO_SIGNED(-191,11),
TO_SIGNED(-236,11),
TO_SIGNED(-280,11),
TO_SIGNED(-323,11),
TO_SIGNED(-365,11),
TO_SIGNED(-406,11),
TO_SIGNED(-444,11),
TO_SIGNED(-481,11),
TO_SIGNED(-516,11),
TO_SIGNED(-549,11),
TO_SIGNED(-580,11),
TO_SIGNED(-609,11),
TO_SIGNED(-635,11),
TO_SIGNED(-659,11),
TO_SIGNED(-680,11),
TO_SIGNED(-699,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-736,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-678,11),
TO_SIGNED(-656,11),
TO_SIGNED(-632,11),
TO_SIGNED(-606,11),
TO_SIGNED(-577,11),
TO_SIGNED(-546,11),
TO_SIGNED(-512,11),
TO_SIGNED(-477,11),
TO_SIGNED(-440,11),
TO_SIGNED(-401,11),
TO_SIGNED(-361,11),
TO_SIGNED(-319,11),
TO_SIGNED(-275,11),
TO_SIGNED(-231,11),
TO_SIGNED(-186,11),
TO_SIGNED(-140,11),
TO_SIGNED(-94,11),
TO_SIGNED(-47,11),
TO_SIGNED(0,11),
TO_SIGNED(47,11),
TO_SIGNED(94,11),
TO_SIGNED(140,11),
TO_SIGNED(186,11),
TO_SIGNED(231,11),
TO_SIGNED(275,11),
TO_SIGNED(319,11),
TO_SIGNED(361,11),
TO_SIGNED(401,11),
TO_SIGNED(440,11),
TO_SIGNED(477,11),
TO_SIGNED(512,11),
TO_SIGNED(546,11),
TO_SIGNED(577,11),
TO_SIGNED(606,11),
TO_SIGNED(632,11),
TO_SIGNED(656,11),
TO_SIGNED(678,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(736,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(699,11),
TO_SIGNED(680,11),
TO_SIGNED(659,11),
TO_SIGNED(635,11),
TO_SIGNED(609,11),
TO_SIGNED(580,11),
TO_SIGNED(549,11),
TO_SIGNED(516,11),
TO_SIGNED(481,11),
TO_SIGNED(444,11),
TO_SIGNED(406,11),
TO_SIGNED(365,11),
TO_SIGNED(323,11),
TO_SIGNED(280,11),
TO_SIGNED(236,11),
TO_SIGNED(191,11),
TO_SIGNED(145,11),
TO_SIGNED(99,11),
TO_SIGNED(52,11),
TO_SIGNED(5,11),
TO_SIGNED(-42,11),
TO_SIGNED(-88,11),
TO_SIGNED(-135,11),
TO_SIGNED(-181,11),
TO_SIGNED(-226,11),
TO_SIGNED(-271,11),
TO_SIGNED(-314,11),
TO_SIGNED(-356,11),
TO_SIGNED(-397,11),
TO_SIGNED(-436,11),
TO_SIGNED(-473,11),
TO_SIGNED(-509,11),
TO_SIGNED(-542,11),
TO_SIGNED(-574,11),
TO_SIGNED(-603,11),
TO_SIGNED(-629,11),
TO_SIGNED(-654,11),
TO_SIGNED(-675,11),
TO_SIGNED(-695,11),
TO_SIGNED(-711,11),
TO_SIGNED(-725,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-716,11),
TO_SIGNED(-700,11),
TO_SIGNED(-682,11),
TO_SIGNED(-661,11),
TO_SIGNED(-638,11),
TO_SIGNED(-612,11),
TO_SIGNED(-584,11),
TO_SIGNED(-553,11),
TO_SIGNED(-520,11),
TO_SIGNED(-485,11),
TO_SIGNED(-449,11),
TO_SIGNED(-410,11),
TO_SIGNED(-370,11),
TO_SIGNED(-328,11),
TO_SIGNED(-285,11),
TO_SIGNED(-241,11),
TO_SIGNED(-196,11),
TO_SIGNED(-151,11),
TO_SIGNED(-104,11),
TO_SIGNED(-58,11),
TO_SIGNED(-11,11),
TO_SIGNED(36,11),
TO_SIGNED(83,11),
TO_SIGNED(130,11),
TO_SIGNED(176,11),
TO_SIGNED(221,11),
TO_SIGNED(266,11),
TO_SIGNED(309,11),
TO_SIGNED(351,11),
TO_SIGNED(392,11),
TO_SIGNED(431,11),
TO_SIGNED(469,11),
TO_SIGNED(505,11),
TO_SIGNED(538,11),
TO_SIGNED(570,11),
TO_SIGNED(599,11),
TO_SIGNED(627,11),
TO_SIGNED(651,11),
TO_SIGNED(673,11),
TO_SIGNED(693,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(739,11),
TO_SIGNED(730,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(685,11),
TO_SIGNED(664,11),
TO_SIGNED(641,11),
TO_SIGNED(615,11),
TO_SIGNED(587,11),
TO_SIGNED(557,11),
TO_SIGNED(524,11),
TO_SIGNED(489,11),
TO_SIGNED(453,11),
TO_SIGNED(415,11),
TO_SIGNED(375,11),
TO_SIGNED(333,11),
TO_SIGNED(290,11),
TO_SIGNED(246,11),
TO_SIGNED(202,11),
TO_SIGNED(156,11),
TO_SIGNED(110,11),
TO_SIGNED(63,11),
TO_SIGNED(16,11),
TO_SIGNED(-31,11),
TO_SIGNED(-78,11),
TO_SIGNED(-124,11),
TO_SIGNED(-171,11),
TO_SIGNED(-216,11),
TO_SIGNED(-261,11),
TO_SIGNED(-304,11),
TO_SIGNED(-346,11),
TO_SIGNED(-387,11),
TO_SIGNED(-427,11),
TO_SIGNED(-465,11),
TO_SIGNED(-501,11),
TO_SIGNED(-535,11),
TO_SIGNED(-567,11),
TO_SIGNED(-596,11),
TO_SIGNED(-624,11),
TO_SIGNED(-648,11),
TO_SIGNED(-671,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-719,11),
TO_SIGNED(-704,11),
TO_SIGNED(-687,11),
TO_SIGNED(-666,11),
TO_SIGNED(-644,11),
TO_SIGNED(-618,11),
TO_SIGNED(-590,11),
TO_SIGNED(-560,11),
TO_SIGNED(-528,11),
TO_SIGNED(-493,11),
TO_SIGNED(-457,11),
TO_SIGNED(-419,11),
TO_SIGNED(-379,11),
TO_SIGNED(-338,11),
TO_SIGNED(-295,11),
TO_SIGNED(-251,11),
TO_SIGNED(-207,11),
TO_SIGNED(-161,11),
TO_SIGNED(-115,11),
TO_SIGNED(-68,11),
TO_SIGNED(-21,11),
TO_SIGNED(26,11),
TO_SIGNED(73,11),
TO_SIGNED(119,11),
TO_SIGNED(165,11),
TO_SIGNED(211,11),
TO_SIGNED(256,11),
TO_SIGNED(299,11),
TO_SIGNED(342,11),
TO_SIGNED(383,11),
TO_SIGNED(422,11),
TO_SIGNED(460,11),
TO_SIGNED(497,11),
TO_SIGNED(531,11),
TO_SIGNED(563,11),
TO_SIGNED(593,11),
TO_SIGNED(621,11),
TO_SIGNED(646,11),
TO_SIGNED(668,11),
TO_SIGNED(688,11),
TO_SIGNED(706,11),
TO_SIGNED(720,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(721,11),
TO_SIGNED(706,11),
TO_SIGNED(689,11),
TO_SIGNED(669,11),
TO_SIGNED(646,11),
TO_SIGNED(621,11),
TO_SIGNED(594,11),
TO_SIGNED(564,11),
TO_SIGNED(532,11),
TO_SIGNED(497,11),
TO_SIGNED(461,11),
TO_SIGNED(423,11),
TO_SIGNED(384,11),
TO_SIGNED(343,11),
TO_SIGNED(300,11),
TO_SIGNED(257,11),
TO_SIGNED(212,11),
TO_SIGNED(166,11),
TO_SIGNED(120,11),
TO_SIGNED(74,11),
TO_SIGNED(27,11),
TO_SIGNED(-20,11),
TO_SIGNED(-67,11),
TO_SIGNED(-114,11),
TO_SIGNED(-160,11),
TO_SIGNED(-206,11),
TO_SIGNED(-250,11),
TO_SIGNED(-294,11),
TO_SIGNED(-337,11),
TO_SIGNED(-378,11),
TO_SIGNED(-418,11),
TO_SIGNED(-456,11),
TO_SIGNED(-493,11),
TO_SIGNED(-527,11),
TO_SIGNED(-559,11),
TO_SIGNED(-590,11),
TO_SIGNED(-618,11),
TO_SIGNED(-643,11),
TO_SIGNED(-666,11),
TO_SIGNED(-686,11),
TO_SIGNED(-704,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-733,11),
TO_SIGNED(-722,11),
TO_SIGNED(-708,11),
TO_SIGNED(-691,11),
TO_SIGNED(-671,11),
TO_SIGNED(-649,11),
TO_SIGNED(-624,11),
TO_SIGNED(-597,11),
TO_SIGNED(-567,11),
TO_SIGNED(-535,11),
TO_SIGNED(-501,11),
TO_SIGNED(-466,11),
TO_SIGNED(-428,11),
TO_SIGNED(-388,11),
TO_SIGNED(-347,11),
TO_SIGNED(-305,11),
TO_SIGNED(-262,11),
TO_SIGNED(-217,11),
TO_SIGNED(-172,11),
TO_SIGNED(-125,11),
TO_SIGNED(-79,11),
TO_SIGNED(-32,11),
TO_SIGNED(15,11),
TO_SIGNED(62,11),
TO_SIGNED(109,11),
TO_SIGNED(155,11),
TO_SIGNED(201,11),
TO_SIGNED(245,11),
TO_SIGNED(289,11),
TO_SIGNED(332,11),
TO_SIGNED(374,11),
TO_SIGNED(414,11),
TO_SIGNED(452,11),
TO_SIGNED(489,11),
TO_SIGNED(523,11),
TO_SIGNED(556,11),
TO_SIGNED(586,11),
TO_SIGNED(615,11),
TO_SIGNED(640,11),
TO_SIGNED(663,11),
TO_SIGNED(684,11),
TO_SIGNED(702,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(710,11),
TO_SIGNED(693,11),
TO_SIGNED(674,11),
TO_SIGNED(652,11),
TO_SIGNED(627,11),
TO_SIGNED(600,11),
TO_SIGNED(571,11),
TO_SIGNED(539,11),
TO_SIGNED(505,11),
TO_SIGNED(470,11),
TO_SIGNED(432,11),
TO_SIGNED(393,11),
TO_SIGNED(352,11),
TO_SIGNED(310,11),
TO_SIGNED(267,11),
TO_SIGNED(222,11),
TO_SIGNED(177,11),
TO_SIGNED(131,11),
TO_SIGNED(84,11),
TO_SIGNED(37,11),
TO_SIGNED(-10,11),
TO_SIGNED(-57,11),
TO_SIGNED(-103,11),
TO_SIGNED(-150,11),
TO_SIGNED(-195,11),
TO_SIGNED(-240,11),
TO_SIGNED(-284,11),
TO_SIGNED(-327,11),
TO_SIGNED(-369,11),
TO_SIGNED(-409,11),
TO_SIGNED(-448,11),
TO_SIGNED(-485,11),
TO_SIGNED(-519,11),
TO_SIGNED(-552,11),
TO_SIGNED(-583,11),
TO_SIGNED(-611,11),
TO_SIGNED(-637,11),
TO_SIGNED(-661,11),
TO_SIGNED(-682,11),
TO_SIGNED(-700,11),
TO_SIGNED(-716,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-725,11),
TO_SIGNED(-711,11),
TO_SIGNED(-695,11),
TO_SIGNED(-676,11),
TO_SIGNED(-654,11),
TO_SIGNED(-630,11),
TO_SIGNED(-603,11),
TO_SIGNED(-574,11),
TO_SIGNED(-543,11),
TO_SIGNED(-509,11),
TO_SIGNED(-474,11),
TO_SIGNED(-437,11),
TO_SIGNED(-397,11),
TO_SIGNED(-357,11),
TO_SIGNED(-315,11),
TO_SIGNED(-272,11),
TO_SIGNED(-227,11),
TO_SIGNED(-182,11),
TO_SIGNED(-136,11),
TO_SIGNED(-90,11),
TO_SIGNED(-43,11),
TO_SIGNED(4,11),
TO_SIGNED(51,11),
TO_SIGNED(98,11),
TO_SIGNED(144,11),
TO_SIGNED(190,11),
TO_SIGNED(235,11),
TO_SIGNED(279,11),
TO_SIGNED(323,11),
TO_SIGNED(364,11),
TO_SIGNED(405,11),
TO_SIGNED(443,11),
TO_SIGNED(480,11),
TO_SIGNED(516,11),
TO_SIGNED(549,11),
TO_SIGNED(580,11),
TO_SIGNED(608,11),
TO_SIGNED(635,11),
TO_SIGNED(658,11),
TO_SIGNED(680,11),
TO_SIGNED(698,11),
TO_SIGNED(714,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(713,11),
TO_SIGNED(697,11),
TO_SIGNED(678,11),
TO_SIGNED(657,11),
TO_SIGNED(633,11),
TO_SIGNED(606,11),
TO_SIGNED(578,11),
TO_SIGNED(547,11),
TO_SIGNED(513,11),
TO_SIGNED(478,11),
TO_SIGNED(441,11),
TO_SIGNED(402,11),
TO_SIGNED(362,11),
TO_SIGNED(320,11),
TO_SIGNED(276,11),
TO_SIGNED(232,11),
TO_SIGNED(187,11),
TO_SIGNED(141,11),
TO_SIGNED(95,11),
TO_SIGNED(48,11),
TO_SIGNED(1,11),
TO_SIGNED(-46,11),
TO_SIGNED(-93,11),
TO_SIGNED(-139,11),
TO_SIGNED(-185,11),
TO_SIGNED(-230,11),
TO_SIGNED(-275,11),
TO_SIGNED(-318,11),
TO_SIGNED(-360,11),
TO_SIGNED(-400,11),
TO_SIGNED(-439,11),
TO_SIGNED(-476,11),
TO_SIGNED(-512,11),
TO_SIGNED(-545,11),
TO_SIGNED(-576,11),
TO_SIGNED(-605,11),
TO_SIGNED(-632,11),
TO_SIGNED(-656,11),
TO_SIGNED(-677,11),
TO_SIGNED(-696,11),
TO_SIGNED(-712,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-715,11),
TO_SIGNED(-699,11),
TO_SIGNED(-681,11),
TO_SIGNED(-659,11),
TO_SIGNED(-636,11),
TO_SIGNED(-610,11),
TO_SIGNED(-581,11),
TO_SIGNED(-550,11),
TO_SIGNED(-517,11),
TO_SIGNED(-482,11),
TO_SIGNED(-445,11),
TO_SIGNED(-406,11),
TO_SIGNED(-366,11),
TO_SIGNED(-324,11),
TO_SIGNED(-281,11),
TO_SIGNED(-237,11),
TO_SIGNED(-192,11),
TO_SIGNED(-147,11),
TO_SIGNED(-100,11),
TO_SIGNED(-53,11),
TO_SIGNED(-6,11),
TO_SIGNED(41,11),
TO_SIGNED(87,11),
TO_SIGNED(134,11),
TO_SIGNED(180,11),
TO_SIGNED(225,11),
TO_SIGNED(270,11),
TO_SIGNED(313,11),
TO_SIGNED(355,11),
TO_SIGNED(396,11),
TO_SIGNED(435,11),
TO_SIGNED(472,11),
TO_SIGNED(508,11),
TO_SIGNED(541,11),
TO_SIGNED(573,11),
TO_SIGNED(602,11),
TO_SIGNED(629,11),
TO_SIGNED(653,11),
TO_SIGNED(675,11),
TO_SIGNED(694,11),
TO_SIGNED(711,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(729,11),
TO_SIGNED(716,11),
TO_SIGNED(701,11),
TO_SIGNED(683,11),
TO_SIGNED(662,11),
TO_SIGNED(639,11),
TO_SIGNED(613,11),
TO_SIGNED(584,11),
TO_SIGNED(554,11),
TO_SIGNED(521,11),
TO_SIGNED(486,11),
TO_SIGNED(449,11),
TO_SIGNED(411,11),
TO_SIGNED(371,11),
TO_SIGNED(329,11),
TO_SIGNED(286,11),
TO_SIGNED(242,11),
TO_SIGNED(197,11),
TO_SIGNED(152,11),
TO_SIGNED(105,11),
TO_SIGNED(59,11),
TO_SIGNED(12,11),
TO_SIGNED(-35,11),
TO_SIGNED(-82,11),
TO_SIGNED(-129,11),
TO_SIGNED(-175,11),
TO_SIGNED(-220,11),
TO_SIGNED(-265,11),
TO_SIGNED(-308,11),
TO_SIGNED(-350,11),
TO_SIGNED(-391,11),
TO_SIGNED(-430,11),
TO_SIGNED(-468,11),
TO_SIGNED(-504,11),
TO_SIGNED(-538,11),
TO_SIGNED(-569,11),
TO_SIGNED(-599,11),
TO_SIGNED(-626,11),
TO_SIGNED(-651,11),
TO_SIGNED(-673,11),
TO_SIGNED(-692,11),
TO_SIGNED(-709,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-685,11),
TO_SIGNED(-664,11),
TO_SIGNED(-641,11),
TO_SIGNED(-616,11),
TO_SIGNED(-588,11),
TO_SIGNED(-557,11),
TO_SIGNED(-525,11),
TO_SIGNED(-490,11),
TO_SIGNED(-454,11),
TO_SIGNED(-415,11),
TO_SIGNED(-375,11),
TO_SIGNED(-334,11),
TO_SIGNED(-291,11),
TO_SIGNED(-247,11),
TO_SIGNED(-203,11),
TO_SIGNED(-157,11),
TO_SIGNED(-111,11),
TO_SIGNED(-64,11),
TO_SIGNED(-17,11),
TO_SIGNED(30,11),
TO_SIGNED(77,11),
TO_SIGNED(123,11),
TO_SIGNED(169,11),
TO_SIGNED(215,11),
TO_SIGNED(260,11),
TO_SIGNED(303,11),
TO_SIGNED(345,11),
TO_SIGNED(387,11),
TO_SIGNED(426,11),
TO_SIGNED(464,11),
TO_SIGNED(500,11),
TO_SIGNED(534,11),
TO_SIGNED(566,11),
TO_SIGNED(596,11),
TO_SIGNED(623,11),
TO_SIGNED(648,11),
TO_SIGNED(670,11),
TO_SIGNED(690,11),
TO_SIGNED(707,11),
TO_SIGNED(721,11),
TO_SIGNED(733,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(705,11),
TO_SIGNED(687,11),
TO_SIGNED(667,11),
TO_SIGNED(644,11),
TO_SIGNED(619,11),
TO_SIGNED(591,11),
TO_SIGNED(561,11),
TO_SIGNED(529,11),
TO_SIGNED(494,11),
TO_SIGNED(458,11),
TO_SIGNED(420,11),
TO_SIGNED(380,11),
TO_SIGNED(339,11),
TO_SIGNED(296,11),
TO_SIGNED(252,11),
TO_SIGNED(208,11),
TO_SIGNED(162,11),
TO_SIGNED(116,11),
TO_SIGNED(69,11),
TO_SIGNED(22,11),
TO_SIGNED(-25,11),
TO_SIGNED(-71,11),
TO_SIGNED(-118,11),
TO_SIGNED(-164,11),
TO_SIGNED(-210,11),
TO_SIGNED(-255,11),
TO_SIGNED(-298,11),
TO_SIGNED(-341,11),
TO_SIGNED(-382,11),
TO_SIGNED(-422,11),
TO_SIGNED(-460,11),
TO_SIGNED(-496,11),
TO_SIGNED(-530,11),
TO_SIGNED(-562,11),
TO_SIGNED(-592,11),
TO_SIGNED(-620,11),
TO_SIGNED(-645,11),
TO_SIGNED(-668,11),
TO_SIGNED(-688,11),
TO_SIGNED(-705,11),
TO_SIGNED(-720,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-721,11),
TO_SIGNED(-706,11),
TO_SIGNED(-689,11),
TO_SIGNED(-669,11),
TO_SIGNED(-647,11),
TO_SIGNED(-622,11),
TO_SIGNED(-594,11),
TO_SIGNED(-564,11),
TO_SIGNED(-532,11),
TO_SIGNED(-498,11),
TO_SIGNED(-462,11),
TO_SIGNED(-424,11),
TO_SIGNED(-385,11),
TO_SIGNED(-344,11),
TO_SIGNED(-301,11),
TO_SIGNED(-258,11),
TO_SIGNED(-213,11),
TO_SIGNED(-167,11),
TO_SIGNED(-121,11),
TO_SIGNED(-75,11),
TO_SIGNED(-28,11),
TO_SIGNED(19,11),
TO_SIGNED(66,11),
TO_SIGNED(113,11),
TO_SIGNED(159,11),
TO_SIGNED(205,11),
TO_SIGNED(249,11),
TO_SIGNED(293,11),
TO_SIGNED(336,11),
TO_SIGNED(377,11),
TO_SIGNED(417,11),
TO_SIGNED(455,11),
TO_SIGNED(492,11),
TO_SIGNED(526,11),
TO_SIGNED(559,11),
TO_SIGNED(589,11),
TO_SIGNED(617,11),
TO_SIGNED(642,11),
TO_SIGNED(665,11),
TO_SIGNED(686,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(708,11),
TO_SIGNED(691,11),
TO_SIGNED(672,11),
TO_SIGNED(650,11),
TO_SIGNED(625,11),
TO_SIGNED(598,11),
TO_SIGNED(568,11),
TO_SIGNED(536,11),
TO_SIGNED(502,11),
TO_SIGNED(466,11),
TO_SIGNED(429,11),
TO_SIGNED(389,11),
TO_SIGNED(348,11),
TO_SIGNED(306,11),
TO_SIGNED(263,11),
TO_SIGNED(218,11),
TO_SIGNED(173,11),
TO_SIGNED(127,11),
TO_SIGNED(80,11),
TO_SIGNED(33,11),
TO_SIGNED(-14,11),
TO_SIGNED(-61,11),
TO_SIGNED(-108,11),
TO_SIGNED(-154,11),
TO_SIGNED(-200,11),
TO_SIGNED(-244,11),
TO_SIGNED(-288,11),
TO_SIGNED(-331,11),
TO_SIGNED(-373,11),
TO_SIGNED(-413,11),
TO_SIGNED(-451,11),
TO_SIGNED(-488,11),
TO_SIGNED(-523,11),
TO_SIGNED(-555,11),
TO_SIGNED(-586,11),
TO_SIGNED(-614,11),
TO_SIGNED(-640,11),
TO_SIGNED(-663,11),
TO_SIGNED(-684,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-729,11),
TO_SIGNED(-739,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-710,11),
TO_SIGNED(-693,11),
TO_SIGNED(-674,11),
TO_SIGNED(-652,11),
TO_SIGNED(-628,11),
TO_SIGNED(-601,11),
TO_SIGNED(-571,11),
TO_SIGNED(-540,11),
TO_SIGNED(-506,11),
TO_SIGNED(-471,11),
TO_SIGNED(-433,11),
TO_SIGNED(-394,11),
TO_SIGNED(-353,11),
TO_SIGNED(-311,11),
TO_SIGNED(-268,11),
TO_SIGNED(-223,11),
TO_SIGNED(-178,11),
TO_SIGNED(-132,11),
TO_SIGNED(-85,11),
TO_SIGNED(-38,11),
TO_SIGNED(9,11),
TO_SIGNED(56,11),
TO_SIGNED(102,11),
TO_SIGNED(149,11),
TO_SIGNED(194,11),
TO_SIGNED(239,11),
TO_SIGNED(283,11),
TO_SIGNED(326,11),
TO_SIGNED(368,11),
TO_SIGNED(408,11),
TO_SIGNED(447,11),
TO_SIGNED(484,11),
TO_SIGNED(519,11),
TO_SIGNED(552,11),
TO_SIGNED(582,11),
TO_SIGNED(611,11),
TO_SIGNED(637,11),
TO_SIGNED(660,11),
TO_SIGNED(681,11),
TO_SIGNED(700,11),
TO_SIGNED(715,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(736,11),
TO_SIGNED(725,11),
TO_SIGNED(712,11),
TO_SIGNED(695,11),
TO_SIGNED(676,11),
TO_SIGNED(655,11),
TO_SIGNED(631,11),
TO_SIGNED(604,11),
TO_SIGNED(575,11),
TO_SIGNED(544,11),
TO_SIGNED(510,11),
TO_SIGNED(475,11),
TO_SIGNED(437,11),
TO_SIGNED(398,11),
TO_SIGNED(358,11),
TO_SIGNED(316,11),
TO_SIGNED(273,11),
TO_SIGNED(228,11),
TO_SIGNED(183,11),
TO_SIGNED(137,11),
TO_SIGNED(91,11),
TO_SIGNED(44,11),
TO_SIGNED(-3,11),
TO_SIGNED(-50,11),
TO_SIGNED(-97,11),
TO_SIGNED(-143,11),
TO_SIGNED(-189,11),
TO_SIGNED(-234,11),
TO_SIGNED(-278,11),
TO_SIGNED(-322,11),
TO_SIGNED(-363,11),
TO_SIGNED(-404,11),
TO_SIGNED(-443,11),
TO_SIGNED(-480,11),
TO_SIGNED(-515,11),
TO_SIGNED(-548,11),
TO_SIGNED(-579,11),
TO_SIGNED(-608,11),
TO_SIGNED(-634,11),
TO_SIGNED(-658,11),
TO_SIGNED(-679,11),
TO_SIGNED(-698,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-679,11),
TO_SIGNED(-657,11),
TO_SIGNED(-633,11),
TO_SIGNED(-607,11),
TO_SIGNED(-578,11),
TO_SIGNED(-547,11),
TO_SIGNED(-514,11),
TO_SIGNED(-479,11),
TO_SIGNED(-442,11),
TO_SIGNED(-403,11),
TO_SIGNED(-362,11),
TO_SIGNED(-321,11),
TO_SIGNED(-277,11),
TO_SIGNED(-233,11),
TO_SIGNED(-188,11),
TO_SIGNED(-142,11),
TO_SIGNED(-96,11),
TO_SIGNED(-49,11),
TO_SIGNED(-2,11),
TO_SIGNED(45,11),
TO_SIGNED(92,11),
TO_SIGNED(138,11),
TO_SIGNED(184,11),
TO_SIGNED(229,11),
TO_SIGNED(274,11),
TO_SIGNED(317,11),
TO_SIGNED(359,11),
TO_SIGNED(399,11),
TO_SIGNED(438,11),
TO_SIGNED(476,11),
TO_SIGNED(511,11),
TO_SIGNED(544,11),
TO_SIGNED(576,11),
TO_SIGNED(605,11),
TO_SIGNED(631,11),
TO_SIGNED(655,11),
TO_SIGNED(677,11),
TO_SIGNED(696,11),
TO_SIGNED(712,11),
TO_SIGNED(725,11),
TO_SIGNED(736,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(715,11),
TO_SIGNED(699,11),
TO_SIGNED(681,11),
TO_SIGNED(660,11),
TO_SIGNED(636,11),
TO_SIGNED(610,11),
TO_SIGNED(582,11),
TO_SIGNED(551,11),
TO_SIGNED(518,11),
TO_SIGNED(483,11),
TO_SIGNED(446,11),
TO_SIGNED(407,11),
TO_SIGNED(367,11),
TO_SIGNED(325,11),
TO_SIGNED(282,11),
TO_SIGNED(238,11),
TO_SIGNED(193,11),
TO_SIGNED(148,11),
TO_SIGNED(101,11),
TO_SIGNED(54,11),
TO_SIGNED(7,11),
TO_SIGNED(-40,11),
TO_SIGNED(-86,11),
TO_SIGNED(-133,11),
TO_SIGNED(-179,11),
TO_SIGNED(-224,11),
TO_SIGNED(-269,11),
TO_SIGNED(-312,11),
TO_SIGNED(-354,11),
TO_SIGNED(-395,11),
TO_SIGNED(-434,11),
TO_SIGNED(-471,11),
TO_SIGNED(-507,11),
TO_SIGNED(-541,11),
TO_SIGNED(-572,11),
TO_SIGNED(-601,11),
TO_SIGNED(-628,11),
TO_SIGNED(-653,11),
TO_SIGNED(-675,11),
TO_SIGNED(-694,11),
TO_SIGNED(-710,11),
TO_SIGNED(-724,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-701,11),
TO_SIGNED(-683,11),
TO_SIGNED(-662,11),
TO_SIGNED(-639,11),
TO_SIGNED(-613,11),
TO_SIGNED(-585,11),
TO_SIGNED(-554,11),
TO_SIGNED(-522,11),
TO_SIGNED(-487,11),
TO_SIGNED(-450,11),
TO_SIGNED(-412,11),
TO_SIGNED(-372,11),
TO_SIGNED(-330,11),
TO_SIGNED(-287,11),
TO_SIGNED(-243,11),
TO_SIGNED(-198,11),
TO_SIGNED(-153,11),
TO_SIGNED(-106,11),
TO_SIGNED(-60,11),
TO_SIGNED(-13,11),
TO_SIGNED(34,11),
TO_SIGNED(81,11),
TO_SIGNED(128,11),
TO_SIGNED(174,11),
TO_SIGNED(219,11),
TO_SIGNED(264,11),
TO_SIGNED(307,11),
TO_SIGNED(349,11),
TO_SIGNED(390,11),
TO_SIGNED(430,11),
TO_SIGNED(467,11),
TO_SIGNED(503,11),
TO_SIGNED(537,11),
TO_SIGNED(569,11),
TO_SIGNED(598,11),
TO_SIGNED(625,11),
TO_SIGNED(650,11),
TO_SIGNED(672,11),
TO_SIGNED(692,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(730,11),
TO_SIGNED(718,11),
TO_SIGNED(703,11),
TO_SIGNED(685,11),
TO_SIGNED(665,11),
TO_SIGNED(642,11),
TO_SIGNED(616,11),
TO_SIGNED(588,11),
TO_SIGNED(558,11),
TO_SIGNED(526,11),
TO_SIGNED(491,11),
TO_SIGNED(455,11),
TO_SIGNED(416,11),
TO_SIGNED(376,11),
TO_SIGNED(335,11),
TO_SIGNED(292,11),
TO_SIGNED(248,11),
TO_SIGNED(204,11),
TO_SIGNED(158,11),
TO_SIGNED(112,11),
TO_SIGNED(65,11),
TO_SIGNED(18,11),
TO_SIGNED(-29,11),
TO_SIGNED(-76,11),
TO_SIGNED(-122,11),
TO_SIGNED(-168,11),
TO_SIGNED(-214,11),
TO_SIGNED(-259,11),
TO_SIGNED(-302,11),
TO_SIGNED(-345,11),
TO_SIGNED(-386,11),
TO_SIGNED(-425,11),
TO_SIGNED(-463,11),
TO_SIGNED(-499,11),
TO_SIGNED(-533,11),
TO_SIGNED(-565,11),
TO_SIGNED(-595,11),
TO_SIGNED(-622,11),
TO_SIGNED(-647,11),
TO_SIGNED(-670,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-721,11),
TO_SIGNED(-733,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-720,11),
TO_SIGNED(-705,11),
TO_SIGNED(-688,11),
TO_SIGNED(-667,11),
TO_SIGNED(-645,11),
TO_SIGNED(-619,11),
TO_SIGNED(-592,11),
TO_SIGNED(-562,11),
TO_SIGNED(-529,11),
TO_SIGNED(-495,11),
TO_SIGNED(-459,11),
TO_SIGNED(-421,11),
TO_SIGNED(-381,11),
TO_SIGNED(-340,11),
TO_SIGNED(-297,11),
TO_SIGNED(-254,11),
TO_SIGNED(-209,11),
TO_SIGNED(-163,11),
TO_SIGNED(-117,11),
TO_SIGNED(-70,11),
TO_SIGNED(-24,11),
TO_SIGNED(24,11),
TO_SIGNED(70,11),
TO_SIGNED(117,11),
TO_SIGNED(163,11),
TO_SIGNED(209,11),
TO_SIGNED(254,11),
TO_SIGNED(297,11),
TO_SIGNED(340,11),
TO_SIGNED(381,11),
TO_SIGNED(421,11),
TO_SIGNED(459,11),
TO_SIGNED(495,11),
TO_SIGNED(529,11),
TO_SIGNED(562,11),
TO_SIGNED(592,11),
TO_SIGNED(619,11),
TO_SIGNED(645,11),
TO_SIGNED(667,11),
TO_SIGNED(688,11),
TO_SIGNED(705,11),
TO_SIGNED(720,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(733,11),
TO_SIGNED(721,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(670,11),
TO_SIGNED(647,11),
TO_SIGNED(622,11),
TO_SIGNED(595,11),
TO_SIGNED(565,11),
TO_SIGNED(533,11),
TO_SIGNED(499,11),
TO_SIGNED(463,11),
TO_SIGNED(425,11),
TO_SIGNED(386,11),
TO_SIGNED(345,11),
TO_SIGNED(302,11),
TO_SIGNED(259,11),
TO_SIGNED(214,11),
TO_SIGNED(168,11),
TO_SIGNED(122,11),
TO_SIGNED(76,11),
TO_SIGNED(29,11),
TO_SIGNED(-18,11),
TO_SIGNED(-65,11),
TO_SIGNED(-112,11),
TO_SIGNED(-158,11),
TO_SIGNED(-204,11),
TO_SIGNED(-248,11),
TO_SIGNED(-292,11),
TO_SIGNED(-335,11),
TO_SIGNED(-376,11),
TO_SIGNED(-416,11),
TO_SIGNED(-455,11),
TO_SIGNED(-491,11),
TO_SIGNED(-526,11),
TO_SIGNED(-558,11),
TO_SIGNED(-588,11),
TO_SIGNED(-616,11),
TO_SIGNED(-642,11),
TO_SIGNED(-665,11),
TO_SIGNED(-685,11),
TO_SIGNED(-703,11),
TO_SIGNED(-718,11),
TO_SIGNED(-730,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-692,11),
TO_SIGNED(-672,11),
TO_SIGNED(-650,11),
TO_SIGNED(-625,11),
TO_SIGNED(-598,11),
TO_SIGNED(-569,11),
TO_SIGNED(-537,11),
TO_SIGNED(-503,11),
TO_SIGNED(-467,11),
TO_SIGNED(-430,11),
TO_SIGNED(-390,11),
TO_SIGNED(-349,11),
TO_SIGNED(-307,11),
TO_SIGNED(-264,11),
TO_SIGNED(-219,11),
TO_SIGNED(-174,11),
TO_SIGNED(-128,11),
TO_SIGNED(-81,11),
TO_SIGNED(-34,11),
TO_SIGNED(13,11),
TO_SIGNED(60,11),
TO_SIGNED(106,11),
TO_SIGNED(153,11),
TO_SIGNED(198,11),
TO_SIGNED(243,11),
TO_SIGNED(287,11),
TO_SIGNED(330,11),
TO_SIGNED(372,11),
TO_SIGNED(412,11),
TO_SIGNED(450,11),
TO_SIGNED(487,11),
TO_SIGNED(522,11),
TO_SIGNED(554,11),
TO_SIGNED(585,11),
TO_SIGNED(613,11),
TO_SIGNED(639,11),
TO_SIGNED(662,11),
TO_SIGNED(683,11),
TO_SIGNED(701,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(724,11),
TO_SIGNED(710,11),
TO_SIGNED(694,11),
TO_SIGNED(675,11),
TO_SIGNED(653,11),
TO_SIGNED(628,11),
TO_SIGNED(601,11),
TO_SIGNED(572,11),
TO_SIGNED(541,11),
TO_SIGNED(507,11),
TO_SIGNED(471,11),
TO_SIGNED(434,11),
TO_SIGNED(395,11),
TO_SIGNED(354,11),
TO_SIGNED(312,11),
TO_SIGNED(269,11),
TO_SIGNED(224,11),
TO_SIGNED(179,11),
TO_SIGNED(133,11),
TO_SIGNED(86,11),
TO_SIGNED(40,11),
TO_SIGNED(-7,11),
TO_SIGNED(-54,11),
TO_SIGNED(-101,11),
TO_SIGNED(-148,11),
TO_SIGNED(-193,11),
TO_SIGNED(-238,11),
TO_SIGNED(-282,11),
TO_SIGNED(-325,11),
TO_SIGNED(-367,11),
TO_SIGNED(-407,11),
TO_SIGNED(-446,11),
TO_SIGNED(-483,11),
TO_SIGNED(-518,11),
TO_SIGNED(-551,11),
TO_SIGNED(-582,11),
TO_SIGNED(-610,11),
TO_SIGNED(-636,11),
TO_SIGNED(-660,11),
TO_SIGNED(-681,11),
TO_SIGNED(-699,11),
TO_SIGNED(-715,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-736,11),
TO_SIGNED(-725,11),
TO_SIGNED(-712,11),
TO_SIGNED(-696,11),
TO_SIGNED(-677,11),
TO_SIGNED(-655,11),
TO_SIGNED(-631,11),
TO_SIGNED(-605,11),
TO_SIGNED(-576,11),
TO_SIGNED(-544,11),
TO_SIGNED(-511,11),
TO_SIGNED(-476,11),
TO_SIGNED(-438,11),
TO_SIGNED(-399,11),
TO_SIGNED(-359,11),
TO_SIGNED(-317,11),
TO_SIGNED(-274,11),
TO_SIGNED(-229,11),
TO_SIGNED(-184,11),
TO_SIGNED(-138,11),
TO_SIGNED(-92,11),
TO_SIGNED(-45,11),
TO_SIGNED(2,11),
TO_SIGNED(49,11),
TO_SIGNED(96,11),
TO_SIGNED(142,11),
TO_SIGNED(188,11),
TO_SIGNED(233,11),
TO_SIGNED(277,11),
TO_SIGNED(321,11),
TO_SIGNED(362,11),
TO_SIGNED(403,11),
TO_SIGNED(442,11),
TO_SIGNED(479,11),
TO_SIGNED(514,11),
TO_SIGNED(547,11),
TO_SIGNED(578,11),
TO_SIGNED(607,11),
TO_SIGNED(633,11),
TO_SIGNED(657,11),
TO_SIGNED(679,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(698,11),
TO_SIGNED(679,11),
TO_SIGNED(658,11),
TO_SIGNED(634,11),
TO_SIGNED(608,11),
TO_SIGNED(579,11),
TO_SIGNED(548,11),
TO_SIGNED(515,11),
TO_SIGNED(480,11),
TO_SIGNED(443,11),
TO_SIGNED(404,11),
TO_SIGNED(363,11),
TO_SIGNED(322,11),
TO_SIGNED(278,11),
TO_SIGNED(234,11),
TO_SIGNED(189,11),
TO_SIGNED(143,11),
TO_SIGNED(97,11),
TO_SIGNED(50,11),
TO_SIGNED(3,11),
TO_SIGNED(-44,11),
TO_SIGNED(-91,11),
TO_SIGNED(-137,11),
TO_SIGNED(-183,11),
TO_SIGNED(-228,11),
TO_SIGNED(-273,11),
TO_SIGNED(-316,11),
TO_SIGNED(-358,11),
TO_SIGNED(-398,11),
TO_SIGNED(-437,11),
TO_SIGNED(-475,11),
TO_SIGNED(-510,11),
TO_SIGNED(-544,11),
TO_SIGNED(-575,11),
TO_SIGNED(-604,11),
TO_SIGNED(-631,11),
TO_SIGNED(-655,11),
TO_SIGNED(-676,11),
TO_SIGNED(-695,11),
TO_SIGNED(-712,11),
TO_SIGNED(-725,11),
TO_SIGNED(-736,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-715,11),
TO_SIGNED(-700,11),
TO_SIGNED(-681,11),
TO_SIGNED(-660,11),
TO_SIGNED(-637,11),
TO_SIGNED(-611,11),
TO_SIGNED(-582,11),
TO_SIGNED(-552,11),
TO_SIGNED(-519,11),
TO_SIGNED(-484,11),
TO_SIGNED(-447,11),
TO_SIGNED(-408,11),
TO_SIGNED(-368,11),
TO_SIGNED(-326,11),
TO_SIGNED(-283,11),
TO_SIGNED(-239,11),
TO_SIGNED(-194,11),
TO_SIGNED(-149,11),
TO_SIGNED(-102,11),
TO_SIGNED(-56,11),
TO_SIGNED(-9,11),
TO_SIGNED(38,11),
TO_SIGNED(85,11),
TO_SIGNED(132,11),
TO_SIGNED(178,11),
TO_SIGNED(223,11),
TO_SIGNED(268,11),
TO_SIGNED(311,11),
TO_SIGNED(353,11),
TO_SIGNED(394,11),
TO_SIGNED(433,11),
TO_SIGNED(471,11),
TO_SIGNED(506,11),
TO_SIGNED(540,11),
TO_SIGNED(571,11),
TO_SIGNED(601,11),
TO_SIGNED(628,11),
TO_SIGNED(652,11),
TO_SIGNED(674,11),
TO_SIGNED(693,11),
TO_SIGNED(710,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(739,11),
TO_SIGNED(729,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(684,11),
TO_SIGNED(663,11),
TO_SIGNED(640,11),
TO_SIGNED(614,11),
TO_SIGNED(586,11),
TO_SIGNED(555,11),
TO_SIGNED(523,11),
TO_SIGNED(488,11),
TO_SIGNED(451,11),
TO_SIGNED(413,11),
TO_SIGNED(373,11),
TO_SIGNED(331,11),
TO_SIGNED(288,11),
TO_SIGNED(244,11),
TO_SIGNED(200,11),
TO_SIGNED(154,11),
TO_SIGNED(108,11),
TO_SIGNED(61,11),
TO_SIGNED(14,11),
TO_SIGNED(-33,11),
TO_SIGNED(-80,11),
TO_SIGNED(-127,11),
TO_SIGNED(-173,11),
TO_SIGNED(-218,11),
TO_SIGNED(-263,11),
TO_SIGNED(-306,11),
TO_SIGNED(-348,11),
TO_SIGNED(-389,11),
TO_SIGNED(-429,11),
TO_SIGNED(-466,11),
TO_SIGNED(-502,11),
TO_SIGNED(-536,11),
TO_SIGNED(-568,11),
TO_SIGNED(-598,11),
TO_SIGNED(-625,11),
TO_SIGNED(-650,11),
TO_SIGNED(-672,11),
TO_SIGNED(-691,11),
TO_SIGNED(-708,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-686,11),
TO_SIGNED(-665,11),
TO_SIGNED(-642,11),
TO_SIGNED(-617,11),
TO_SIGNED(-589,11),
TO_SIGNED(-559,11),
TO_SIGNED(-526,11),
TO_SIGNED(-492,11),
TO_SIGNED(-455,11),
TO_SIGNED(-417,11),
TO_SIGNED(-377,11),
TO_SIGNED(-336,11),
TO_SIGNED(-293,11),
TO_SIGNED(-249,11),
TO_SIGNED(-205,11),
TO_SIGNED(-159,11),
TO_SIGNED(-113,11),
TO_SIGNED(-66,11),
TO_SIGNED(-19,11),
TO_SIGNED(28,11),
TO_SIGNED(75,11),
TO_SIGNED(121,11),
TO_SIGNED(167,11),
TO_SIGNED(213,11),
TO_SIGNED(258,11),
TO_SIGNED(301,11),
TO_SIGNED(344,11),
TO_SIGNED(385,11),
TO_SIGNED(424,11),
TO_SIGNED(462,11),
TO_SIGNED(498,11),
TO_SIGNED(532,11),
TO_SIGNED(564,11),
TO_SIGNED(594,11),
TO_SIGNED(622,11),
TO_SIGNED(647,11),
TO_SIGNED(669,11),
TO_SIGNED(689,11),
TO_SIGNED(706,11),
TO_SIGNED(721,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(720,11),
TO_SIGNED(705,11),
TO_SIGNED(688,11),
TO_SIGNED(668,11),
TO_SIGNED(645,11),
TO_SIGNED(620,11),
TO_SIGNED(592,11),
TO_SIGNED(562,11),
TO_SIGNED(530,11),
TO_SIGNED(496,11),
TO_SIGNED(460,11),
TO_SIGNED(422,11),
TO_SIGNED(382,11),
TO_SIGNED(341,11),
TO_SIGNED(298,11),
TO_SIGNED(255,11),
TO_SIGNED(210,11),
TO_SIGNED(164,11),
TO_SIGNED(118,11),
TO_SIGNED(71,11),
TO_SIGNED(25,11),
TO_SIGNED(-22,11),
TO_SIGNED(-69,11),
TO_SIGNED(-116,11),
TO_SIGNED(-162,11),
TO_SIGNED(-208,11),
TO_SIGNED(-252,11),
TO_SIGNED(-296,11),
TO_SIGNED(-339,11),
TO_SIGNED(-380,11),
TO_SIGNED(-420,11),
TO_SIGNED(-458,11),
TO_SIGNED(-494,11),
TO_SIGNED(-529,11),
TO_SIGNED(-561,11),
TO_SIGNED(-591,11),
TO_SIGNED(-619,11),
TO_SIGNED(-644,11),
TO_SIGNED(-667,11),
TO_SIGNED(-687,11),
TO_SIGNED(-705,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-733,11),
TO_SIGNED(-721,11),
TO_SIGNED(-707,11),
TO_SIGNED(-690,11),
TO_SIGNED(-670,11),
TO_SIGNED(-648,11),
TO_SIGNED(-623,11),
TO_SIGNED(-596,11),
TO_SIGNED(-566,11),
TO_SIGNED(-534,11),
TO_SIGNED(-500,11),
TO_SIGNED(-464,11),
TO_SIGNED(-426,11),
TO_SIGNED(-387,11),
TO_SIGNED(-345,11),
TO_SIGNED(-303,11),
TO_SIGNED(-260,11),
TO_SIGNED(-215,11),
TO_SIGNED(-169,11),
TO_SIGNED(-123,11),
TO_SIGNED(-77,11),
TO_SIGNED(-30,11),
TO_SIGNED(17,11),
TO_SIGNED(64,11),
TO_SIGNED(111,11),
TO_SIGNED(157,11),
TO_SIGNED(203,11),
TO_SIGNED(247,11),
TO_SIGNED(291,11),
TO_SIGNED(334,11),
TO_SIGNED(375,11),
TO_SIGNED(415,11),
TO_SIGNED(454,11),
TO_SIGNED(490,11),
TO_SIGNED(525,11),
TO_SIGNED(557,11),
TO_SIGNED(588,11),
TO_SIGNED(616,11),
TO_SIGNED(641,11),
TO_SIGNED(664,11),
TO_SIGNED(685,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(709,11),
TO_SIGNED(692,11),
TO_SIGNED(673,11),
TO_SIGNED(651,11),
TO_SIGNED(626,11),
TO_SIGNED(599,11),
TO_SIGNED(569,11),
TO_SIGNED(538,11),
TO_SIGNED(504,11),
TO_SIGNED(468,11),
TO_SIGNED(430,11),
TO_SIGNED(391,11),
TO_SIGNED(350,11),
TO_SIGNED(308,11),
TO_SIGNED(265,11),
TO_SIGNED(220,11),
TO_SIGNED(175,11),
TO_SIGNED(129,11),
TO_SIGNED(82,11),
TO_SIGNED(35,11),
TO_SIGNED(-12,11),
TO_SIGNED(-59,11),
TO_SIGNED(-105,11),
TO_SIGNED(-152,11),
TO_SIGNED(-197,11),
TO_SIGNED(-242,11),
TO_SIGNED(-286,11),
TO_SIGNED(-329,11),
TO_SIGNED(-371,11),
TO_SIGNED(-411,11),
TO_SIGNED(-449,11),
TO_SIGNED(-486,11),
TO_SIGNED(-521,11),
TO_SIGNED(-554,11),
TO_SIGNED(-584,11),
TO_SIGNED(-613,11),
TO_SIGNED(-639,11),
TO_SIGNED(-662,11),
TO_SIGNED(-683,11),
TO_SIGNED(-701,11),
TO_SIGNED(-716,11),
TO_SIGNED(-729,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-711,11),
TO_SIGNED(-694,11),
TO_SIGNED(-675,11),
TO_SIGNED(-653,11),
TO_SIGNED(-629,11),
TO_SIGNED(-602,11),
TO_SIGNED(-573,11),
TO_SIGNED(-541,11),
TO_SIGNED(-508,11),
TO_SIGNED(-472,11),
TO_SIGNED(-435,11),
TO_SIGNED(-396,11),
TO_SIGNED(-355,11),
TO_SIGNED(-313,11),
TO_SIGNED(-270,11),
TO_SIGNED(-225,11),
TO_SIGNED(-180,11),
TO_SIGNED(-134,11),
TO_SIGNED(-87,11),
TO_SIGNED(-41,11),
TO_SIGNED(6,11),
TO_SIGNED(53,11),
TO_SIGNED(100,11),
TO_SIGNED(147,11),
TO_SIGNED(192,11),
TO_SIGNED(237,11),
TO_SIGNED(281,11),
TO_SIGNED(324,11),
TO_SIGNED(366,11),
TO_SIGNED(406,11),
TO_SIGNED(445,11),
TO_SIGNED(482,11),
TO_SIGNED(517,11),
TO_SIGNED(550,11),
TO_SIGNED(581,11),
TO_SIGNED(610,11),
TO_SIGNED(636,11),
TO_SIGNED(659,11),
TO_SIGNED(681,11),
TO_SIGNED(699,11),
TO_SIGNED(715,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(712,11),
TO_SIGNED(696,11),
TO_SIGNED(677,11),
TO_SIGNED(656,11),
TO_SIGNED(632,11),
TO_SIGNED(605,11),
TO_SIGNED(576,11),
TO_SIGNED(545,11),
TO_SIGNED(512,11),
TO_SIGNED(476,11),
TO_SIGNED(439,11),
TO_SIGNED(400,11),
TO_SIGNED(360,11),
TO_SIGNED(318,11),
TO_SIGNED(275,11),
TO_SIGNED(230,11),
TO_SIGNED(185,11),
TO_SIGNED(139,11),
TO_SIGNED(93,11),
TO_SIGNED(46,11),
TO_SIGNED(-1,11),
TO_SIGNED(-48,11),
TO_SIGNED(-95,11),
TO_SIGNED(-141,11),
TO_SIGNED(-187,11),
TO_SIGNED(-232,11),
TO_SIGNED(-276,11),
TO_SIGNED(-320,11),
TO_SIGNED(-362,11),
TO_SIGNED(-402,11),
TO_SIGNED(-441,11),
TO_SIGNED(-478,11),
TO_SIGNED(-513,11),
TO_SIGNED(-547,11),
TO_SIGNED(-578,11),
TO_SIGNED(-606,11),
TO_SIGNED(-633,11),
TO_SIGNED(-657,11),
TO_SIGNED(-678,11),
TO_SIGNED(-697,11),
TO_SIGNED(-713,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-714,11),
TO_SIGNED(-698,11),
TO_SIGNED(-680,11),
TO_SIGNED(-658,11),
TO_SIGNED(-635,11),
TO_SIGNED(-608,11),
TO_SIGNED(-580,11),
TO_SIGNED(-549,11),
TO_SIGNED(-516,11),
TO_SIGNED(-480,11),
TO_SIGNED(-443,11),
TO_SIGNED(-405,11),
TO_SIGNED(-364,11),
TO_SIGNED(-323,11),
TO_SIGNED(-279,11),
TO_SIGNED(-235,11),
TO_SIGNED(-190,11),
TO_SIGNED(-144,11),
TO_SIGNED(-98,11),
TO_SIGNED(-51,11),
TO_SIGNED(-4,11),
TO_SIGNED(43,11),
TO_SIGNED(90,11),
TO_SIGNED(136,11),
TO_SIGNED(182,11),
TO_SIGNED(227,11),
TO_SIGNED(272,11),
TO_SIGNED(315,11),
TO_SIGNED(357,11),
TO_SIGNED(397,11),
TO_SIGNED(437,11),
TO_SIGNED(474,11),
TO_SIGNED(509,11),
TO_SIGNED(543,11),
TO_SIGNED(574,11),
TO_SIGNED(603,11),
TO_SIGNED(630,11),
TO_SIGNED(654,11),
TO_SIGNED(676,11),
TO_SIGNED(695,11),
TO_SIGNED(711,11),
TO_SIGNED(725,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(716,11),
TO_SIGNED(700,11),
TO_SIGNED(682,11),
TO_SIGNED(661,11),
TO_SIGNED(637,11),
TO_SIGNED(611,11),
TO_SIGNED(583,11),
TO_SIGNED(552,11),
TO_SIGNED(519,11),
TO_SIGNED(485,11),
TO_SIGNED(448,11),
TO_SIGNED(409,11),
TO_SIGNED(369,11),
TO_SIGNED(327,11),
TO_SIGNED(284,11),
TO_SIGNED(240,11),
TO_SIGNED(195,11),
TO_SIGNED(150,11),
TO_SIGNED(103,11),
TO_SIGNED(57,11),
TO_SIGNED(10,11),
TO_SIGNED(-37,11),
TO_SIGNED(-84,11),
TO_SIGNED(-131,11),
TO_SIGNED(-177,11),
TO_SIGNED(-222,11),
TO_SIGNED(-267,11),
TO_SIGNED(-310,11),
TO_SIGNED(-352,11),
TO_SIGNED(-393,11),
TO_SIGNED(-432,11),
TO_SIGNED(-470,11),
TO_SIGNED(-505,11),
TO_SIGNED(-539,11),
TO_SIGNED(-571,11),
TO_SIGNED(-600,11),
TO_SIGNED(-627,11),
TO_SIGNED(-652,11),
TO_SIGNED(-674,11),
TO_SIGNED(-693,11),
TO_SIGNED(-710,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-702,11),
TO_SIGNED(-684,11),
TO_SIGNED(-663,11),
TO_SIGNED(-640,11),
TO_SIGNED(-615,11),
TO_SIGNED(-586,11),
TO_SIGNED(-556,11),
TO_SIGNED(-523,11),
TO_SIGNED(-489,11),
TO_SIGNED(-452,11),
TO_SIGNED(-414,11),
TO_SIGNED(-374,11),
TO_SIGNED(-332,11),
TO_SIGNED(-289,11),
TO_SIGNED(-245,11),
TO_SIGNED(-201,11),
TO_SIGNED(-155,11),
TO_SIGNED(-109,11),
TO_SIGNED(-62,11),
TO_SIGNED(-15,11),
TO_SIGNED(32,11),
TO_SIGNED(79,11),
TO_SIGNED(125,11),
TO_SIGNED(172,11),
TO_SIGNED(217,11),
TO_SIGNED(262,11),
TO_SIGNED(305,11),
TO_SIGNED(347,11),
TO_SIGNED(388,11),
TO_SIGNED(428,11),
TO_SIGNED(466,11),
TO_SIGNED(501,11),
TO_SIGNED(535,11),
TO_SIGNED(567,11),
TO_SIGNED(597,11),
TO_SIGNED(624,11),
TO_SIGNED(649,11),
TO_SIGNED(671,11),
TO_SIGNED(691,11),
TO_SIGNED(708,11),
TO_SIGNED(722,11),
TO_SIGNED(733,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(704,11),
TO_SIGNED(686,11),
TO_SIGNED(666,11),
TO_SIGNED(643,11),
TO_SIGNED(618,11),
TO_SIGNED(590,11),
TO_SIGNED(559,11),
TO_SIGNED(527,11),
TO_SIGNED(493,11),
TO_SIGNED(456,11),
TO_SIGNED(418,11),
TO_SIGNED(378,11),
TO_SIGNED(337,11),
TO_SIGNED(294,11),
TO_SIGNED(250,11),
TO_SIGNED(206,11),
TO_SIGNED(160,11),
TO_SIGNED(114,11),
TO_SIGNED(67,11),
TO_SIGNED(20,11),
TO_SIGNED(-27,11),
TO_SIGNED(-74,11),
TO_SIGNED(-120,11),
TO_SIGNED(-166,11),
TO_SIGNED(-212,11),
TO_SIGNED(-257,11),
TO_SIGNED(-300,11),
TO_SIGNED(-343,11),
TO_SIGNED(-384,11),
TO_SIGNED(-423,11),
TO_SIGNED(-461,11),
TO_SIGNED(-497,11),
TO_SIGNED(-532,11),
TO_SIGNED(-564,11),
TO_SIGNED(-594,11),
TO_SIGNED(-621,11),
TO_SIGNED(-646,11),
TO_SIGNED(-669,11),
TO_SIGNED(-689,11),
TO_SIGNED(-706,11),
TO_SIGNED(-721,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-720,11),
TO_SIGNED(-706,11),
TO_SIGNED(-688,11),
TO_SIGNED(-668,11),
TO_SIGNED(-646,11),
TO_SIGNED(-621,11),
TO_SIGNED(-593,11),
TO_SIGNED(-563,11),
TO_SIGNED(-531,11),
TO_SIGNED(-497,11),
TO_SIGNED(-460,11),
TO_SIGNED(-422,11),
TO_SIGNED(-383,11),
TO_SIGNED(-342,11),
TO_SIGNED(-299,11),
TO_SIGNED(-256,11),
TO_SIGNED(-211,11),
TO_SIGNED(-165,11),
TO_SIGNED(-119,11),
TO_SIGNED(-73,11),
TO_SIGNED(-26,11),
TO_SIGNED(21,11),
TO_SIGNED(68,11),
TO_SIGNED(115,11),
TO_SIGNED(161,11),
TO_SIGNED(207,11),
TO_SIGNED(251,11),
TO_SIGNED(295,11),
TO_SIGNED(338,11),
TO_SIGNED(379,11),
TO_SIGNED(419,11),
TO_SIGNED(457,11),
TO_SIGNED(493,11),
TO_SIGNED(528,11),
TO_SIGNED(560,11),
TO_SIGNED(590,11),
TO_SIGNED(618,11),
TO_SIGNED(644,11),
TO_SIGNED(666,11),
TO_SIGNED(687,11),
TO_SIGNED(704,11),
TO_SIGNED(719,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(671,11),
TO_SIGNED(648,11),
TO_SIGNED(624,11),
TO_SIGNED(596,11),
TO_SIGNED(567,11),
TO_SIGNED(535,11),
TO_SIGNED(501,11),
TO_SIGNED(465,11),
TO_SIGNED(427,11),
TO_SIGNED(387,11),
TO_SIGNED(346,11),
TO_SIGNED(304,11),
TO_SIGNED(261,11),
TO_SIGNED(216,11),
TO_SIGNED(171,11),
TO_SIGNED(124,11),
TO_SIGNED(78,11),
TO_SIGNED(31,11),
TO_SIGNED(-16,11),
TO_SIGNED(-63,11),
TO_SIGNED(-110,11),
TO_SIGNED(-156,11),
TO_SIGNED(-202,11),
TO_SIGNED(-246,11),
TO_SIGNED(-290,11),
TO_SIGNED(-333,11),
TO_SIGNED(-375,11),
TO_SIGNED(-415,11),
TO_SIGNED(-453,11),
TO_SIGNED(-489,11),
TO_SIGNED(-524,11),
TO_SIGNED(-557,11),
TO_SIGNED(-587,11),
TO_SIGNED(-615,11),
TO_SIGNED(-641,11),
TO_SIGNED(-664,11),
TO_SIGNED(-685,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-730,11),
TO_SIGNED(-739,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-693,11),
TO_SIGNED(-673,11),
TO_SIGNED(-651,11),
TO_SIGNED(-627,11),
TO_SIGNED(-599,11),
TO_SIGNED(-570,11),
TO_SIGNED(-538,11),
TO_SIGNED(-505,11),
TO_SIGNED(-469,11),
TO_SIGNED(-431,11),
TO_SIGNED(-392,11),
TO_SIGNED(-351,11),
TO_SIGNED(-309,11),
TO_SIGNED(-266,11),
TO_SIGNED(-221,11),
TO_SIGNED(-176,11),
TO_SIGNED(-130,11),
TO_SIGNED(-83,11),
TO_SIGNED(-36,11),
TO_SIGNED(11,11),
TO_SIGNED(58,11),
TO_SIGNED(104,11),
TO_SIGNED(151,11),
TO_SIGNED(196,11),
TO_SIGNED(241,11),
TO_SIGNED(285,11),
TO_SIGNED(328,11),
TO_SIGNED(370,11),
TO_SIGNED(410,11),
TO_SIGNED(449,11),
TO_SIGNED(485,11),
TO_SIGNED(520,11),
TO_SIGNED(553,11),
TO_SIGNED(584,11),
TO_SIGNED(612,11),
TO_SIGNED(638,11),
TO_SIGNED(661,11),
TO_SIGNED(682,11),
TO_SIGNED(700,11),
TO_SIGNED(716,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(725,11),
TO_SIGNED(711,11),
TO_SIGNED(695,11),
TO_SIGNED(675,11),
TO_SIGNED(654,11),
TO_SIGNED(629,11),
TO_SIGNED(603,11),
TO_SIGNED(574,11),
TO_SIGNED(542,11),
TO_SIGNED(509,11),
TO_SIGNED(473,11),
TO_SIGNED(436,11),
TO_SIGNED(397,11),
TO_SIGNED(356,11),
TO_SIGNED(314,11),
TO_SIGNED(271,11),
TO_SIGNED(226,11),
TO_SIGNED(181,11),
TO_SIGNED(135,11),
TO_SIGNED(88,11),
TO_SIGNED(42,11),
TO_SIGNED(-5,11),
TO_SIGNED(-52,11),
TO_SIGNED(-99,11),
TO_SIGNED(-145,11),
TO_SIGNED(-191,11),
TO_SIGNED(-236,11),
TO_SIGNED(-280,11),
TO_SIGNED(-323,11),
TO_SIGNED(-365,11),
TO_SIGNED(-406,11),
TO_SIGNED(-444,11),
TO_SIGNED(-481,11),
TO_SIGNED(-516,11),
TO_SIGNED(-549,11),
TO_SIGNED(-580,11),
TO_SIGNED(-609,11),
TO_SIGNED(-635,11),
TO_SIGNED(-659,11),
TO_SIGNED(-680,11),
TO_SIGNED(-699,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-736,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-678,11),
TO_SIGNED(-656,11),
TO_SIGNED(-632,11),
TO_SIGNED(-606,11),
TO_SIGNED(-577,11),
TO_SIGNED(-546,11),
TO_SIGNED(-512,11),
TO_SIGNED(-477,11),
TO_SIGNED(-440,11),
TO_SIGNED(-401,11),
TO_SIGNED(-361,11),
TO_SIGNED(-319,11),
TO_SIGNED(-275,11),
TO_SIGNED(-231,11),
TO_SIGNED(-186,11),
TO_SIGNED(-140,11),
TO_SIGNED(-94,11),
TO_SIGNED(-47,11),
TO_SIGNED(0,11),
TO_SIGNED(47,11),
TO_SIGNED(94,11),
TO_SIGNED(140,11),
TO_SIGNED(186,11),
TO_SIGNED(231,11),
TO_SIGNED(275,11),
TO_SIGNED(319,11),
TO_SIGNED(361,11),
TO_SIGNED(401,11),
TO_SIGNED(440,11),
TO_SIGNED(477,11),
TO_SIGNED(512,11),
TO_SIGNED(546,11),
TO_SIGNED(577,11),
TO_SIGNED(606,11),
TO_SIGNED(632,11),
TO_SIGNED(656,11),
TO_SIGNED(678,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(736,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(699,11),
TO_SIGNED(680,11),
TO_SIGNED(659,11),
TO_SIGNED(635,11),
TO_SIGNED(609,11),
TO_SIGNED(580,11),
TO_SIGNED(549,11),
TO_SIGNED(516,11),
TO_SIGNED(481,11),
TO_SIGNED(444,11),
TO_SIGNED(406,11),
TO_SIGNED(365,11),
TO_SIGNED(323,11),
TO_SIGNED(280,11),
TO_SIGNED(236,11),
TO_SIGNED(191,11),
TO_SIGNED(145,11),
TO_SIGNED(99,11),
TO_SIGNED(52,11),
TO_SIGNED(5,11),
TO_SIGNED(-42,11),
TO_SIGNED(-88,11),
TO_SIGNED(-135,11),
TO_SIGNED(-181,11),
TO_SIGNED(-226,11),
TO_SIGNED(-271,11),
TO_SIGNED(-314,11),
TO_SIGNED(-356,11),
TO_SIGNED(-397,11),
TO_SIGNED(-436,11),
TO_SIGNED(-473,11),
TO_SIGNED(-509,11),
TO_SIGNED(-542,11),
TO_SIGNED(-574,11),
TO_SIGNED(-603,11),
TO_SIGNED(-629,11),
TO_SIGNED(-654,11),
TO_SIGNED(-675,11),
TO_SIGNED(-695,11),
TO_SIGNED(-711,11),
TO_SIGNED(-725,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-716,11),
TO_SIGNED(-700,11),
TO_SIGNED(-682,11),
TO_SIGNED(-661,11),
TO_SIGNED(-638,11),
TO_SIGNED(-612,11),
TO_SIGNED(-584,11),
TO_SIGNED(-553,11),
TO_SIGNED(-520,11),
TO_SIGNED(-485,11),
TO_SIGNED(-449,11),
TO_SIGNED(-410,11),
TO_SIGNED(-370,11),
TO_SIGNED(-328,11),
TO_SIGNED(-285,11),
TO_SIGNED(-241,11),
TO_SIGNED(-196,11),
TO_SIGNED(-151,11),
TO_SIGNED(-104,11),
TO_SIGNED(-58,11),
TO_SIGNED(-11,11),
TO_SIGNED(36,11),
TO_SIGNED(83,11),
TO_SIGNED(130,11),
TO_SIGNED(176,11),
TO_SIGNED(221,11),
TO_SIGNED(266,11),
TO_SIGNED(309,11),
TO_SIGNED(351,11),
TO_SIGNED(392,11),
TO_SIGNED(431,11),
TO_SIGNED(469,11),
TO_SIGNED(505,11),
TO_SIGNED(538,11),
TO_SIGNED(570,11),
TO_SIGNED(599,11),
TO_SIGNED(627,11),
TO_SIGNED(651,11),
TO_SIGNED(673,11),
TO_SIGNED(693,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(739,11),
TO_SIGNED(730,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(685,11),
TO_SIGNED(664,11),
TO_SIGNED(641,11),
TO_SIGNED(615,11),
TO_SIGNED(587,11),
TO_SIGNED(557,11),
TO_SIGNED(524,11),
TO_SIGNED(489,11),
TO_SIGNED(453,11),
TO_SIGNED(415,11),
TO_SIGNED(375,11),
TO_SIGNED(333,11),
TO_SIGNED(290,11),
TO_SIGNED(246,11),
TO_SIGNED(202,11),
TO_SIGNED(156,11),
TO_SIGNED(110,11),
TO_SIGNED(63,11),
TO_SIGNED(16,11),
TO_SIGNED(-31,11),
TO_SIGNED(-78,11),
TO_SIGNED(-124,11),
TO_SIGNED(-171,11),
TO_SIGNED(-216,11),
TO_SIGNED(-261,11),
TO_SIGNED(-304,11),
TO_SIGNED(-346,11),
TO_SIGNED(-387,11),
TO_SIGNED(-427,11),
TO_SIGNED(-465,11),
TO_SIGNED(-501,11),
TO_SIGNED(-535,11),
TO_SIGNED(-567,11),
TO_SIGNED(-596,11),
TO_SIGNED(-624,11),
TO_SIGNED(-648,11),
TO_SIGNED(-671,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-719,11),
TO_SIGNED(-704,11),
TO_SIGNED(-687,11),
TO_SIGNED(-666,11),
TO_SIGNED(-644,11),
TO_SIGNED(-618,11),
TO_SIGNED(-590,11),
TO_SIGNED(-560,11),
TO_SIGNED(-528,11),
TO_SIGNED(-493,11),
TO_SIGNED(-457,11),
TO_SIGNED(-419,11),
TO_SIGNED(-379,11),
TO_SIGNED(-338,11),
TO_SIGNED(-295,11),
TO_SIGNED(-251,11),
TO_SIGNED(-207,11),
TO_SIGNED(-161,11),
TO_SIGNED(-115,11),
TO_SIGNED(-68,11),
TO_SIGNED(-21,11),
TO_SIGNED(26,11),
TO_SIGNED(73,11),
TO_SIGNED(119,11),
TO_SIGNED(165,11),
TO_SIGNED(211,11),
TO_SIGNED(256,11),
TO_SIGNED(299,11),
TO_SIGNED(342,11),
TO_SIGNED(383,11),
TO_SIGNED(422,11),
TO_SIGNED(460,11),
TO_SIGNED(497,11),
TO_SIGNED(531,11),
TO_SIGNED(563,11),
TO_SIGNED(593,11),
TO_SIGNED(621,11),
TO_SIGNED(646,11),
TO_SIGNED(668,11),
TO_SIGNED(688,11),
TO_SIGNED(706,11),
TO_SIGNED(720,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(721,11),
TO_SIGNED(706,11),
TO_SIGNED(689,11),
TO_SIGNED(669,11),
TO_SIGNED(646,11),
TO_SIGNED(621,11),
TO_SIGNED(594,11),
TO_SIGNED(564,11),
TO_SIGNED(532,11),
TO_SIGNED(497,11),
TO_SIGNED(461,11),
TO_SIGNED(423,11),
TO_SIGNED(384,11),
TO_SIGNED(343,11),
TO_SIGNED(300,11),
TO_SIGNED(257,11),
TO_SIGNED(212,11),
TO_SIGNED(166,11),
TO_SIGNED(120,11),
TO_SIGNED(74,11),
TO_SIGNED(27,11),
TO_SIGNED(-20,11),
TO_SIGNED(-67,11),
TO_SIGNED(-114,11),
TO_SIGNED(-160,11),
TO_SIGNED(-206,11),
TO_SIGNED(-250,11),
TO_SIGNED(-294,11),
TO_SIGNED(-337,11),
TO_SIGNED(-378,11),
TO_SIGNED(-418,11),
TO_SIGNED(-456,11),
TO_SIGNED(-493,11),
TO_SIGNED(-527,11),
TO_SIGNED(-559,11),
TO_SIGNED(-590,11),
TO_SIGNED(-618,11),
TO_SIGNED(-643,11),
TO_SIGNED(-666,11),
TO_SIGNED(-686,11),
TO_SIGNED(-704,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-733,11),
TO_SIGNED(-722,11),
TO_SIGNED(-708,11),
TO_SIGNED(-691,11),
TO_SIGNED(-671,11),
TO_SIGNED(-649,11),
TO_SIGNED(-624,11),
TO_SIGNED(-597,11),
TO_SIGNED(-567,11),
TO_SIGNED(-535,11),
TO_SIGNED(-501,11),
TO_SIGNED(-466,11),
TO_SIGNED(-428,11),
TO_SIGNED(-388,11),
TO_SIGNED(-347,11),
TO_SIGNED(-305,11),
TO_SIGNED(-262,11),
TO_SIGNED(-217,11),
TO_SIGNED(-172,11),
TO_SIGNED(-125,11),
TO_SIGNED(-79,11),
TO_SIGNED(-32,11),
TO_SIGNED(15,11),
TO_SIGNED(62,11),
TO_SIGNED(109,11),
TO_SIGNED(155,11),
TO_SIGNED(201,11),
TO_SIGNED(245,11),
TO_SIGNED(289,11),
TO_SIGNED(332,11),
TO_SIGNED(374,11),
TO_SIGNED(414,11),
TO_SIGNED(452,11),
TO_SIGNED(489,11),
TO_SIGNED(523,11),
TO_SIGNED(556,11),
TO_SIGNED(586,11),
TO_SIGNED(615,11),
TO_SIGNED(640,11),
TO_SIGNED(663,11),
TO_SIGNED(684,11),
TO_SIGNED(702,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(710,11),
TO_SIGNED(693,11),
TO_SIGNED(674,11),
TO_SIGNED(652,11),
TO_SIGNED(627,11),
TO_SIGNED(600,11),
TO_SIGNED(571,11),
TO_SIGNED(539,11),
TO_SIGNED(505,11),
TO_SIGNED(470,11),
TO_SIGNED(432,11),
TO_SIGNED(393,11),
TO_SIGNED(352,11),
TO_SIGNED(310,11),
TO_SIGNED(267,11),
TO_SIGNED(222,11),
TO_SIGNED(177,11),
TO_SIGNED(131,11),
TO_SIGNED(84,11),
TO_SIGNED(37,11),
TO_SIGNED(-10,11),
TO_SIGNED(-57,11),
TO_SIGNED(-103,11),
TO_SIGNED(-150,11),
TO_SIGNED(-195,11),
TO_SIGNED(-240,11),
TO_SIGNED(-284,11),
TO_SIGNED(-327,11),
TO_SIGNED(-369,11),
TO_SIGNED(-409,11),
TO_SIGNED(-448,11),
TO_SIGNED(-485,11),
TO_SIGNED(-519,11),
TO_SIGNED(-552,11),
TO_SIGNED(-583,11),
TO_SIGNED(-611,11),
TO_SIGNED(-637,11),
TO_SIGNED(-661,11),
TO_SIGNED(-682,11),
TO_SIGNED(-700,11),
TO_SIGNED(-716,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-725,11),
TO_SIGNED(-711,11),
TO_SIGNED(-695,11),
TO_SIGNED(-676,11),
TO_SIGNED(-654,11),
TO_SIGNED(-630,11),
TO_SIGNED(-603,11),
TO_SIGNED(-574,11),
TO_SIGNED(-543,11),
TO_SIGNED(-509,11),
TO_SIGNED(-474,11),
TO_SIGNED(-437,11),
TO_SIGNED(-397,11),
TO_SIGNED(-357,11),
TO_SIGNED(-315,11),
TO_SIGNED(-272,11),
TO_SIGNED(-227,11),
TO_SIGNED(-182,11),
TO_SIGNED(-136,11),
TO_SIGNED(-90,11),
TO_SIGNED(-43,11),
TO_SIGNED(4,11),
TO_SIGNED(51,11),
TO_SIGNED(98,11),
TO_SIGNED(144,11),
TO_SIGNED(190,11),
TO_SIGNED(235,11),
TO_SIGNED(279,11),
TO_SIGNED(323,11),
TO_SIGNED(364,11),
TO_SIGNED(405,11),
TO_SIGNED(443,11),
TO_SIGNED(480,11),
TO_SIGNED(516,11),
TO_SIGNED(549,11),
TO_SIGNED(580,11),
TO_SIGNED(608,11),
TO_SIGNED(635,11),
TO_SIGNED(658,11),
TO_SIGNED(680,11),
TO_SIGNED(698,11),
TO_SIGNED(714,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(713,11),
TO_SIGNED(697,11),
TO_SIGNED(678,11),
TO_SIGNED(657,11),
TO_SIGNED(633,11),
TO_SIGNED(606,11),
TO_SIGNED(578,11),
TO_SIGNED(547,11),
TO_SIGNED(513,11),
TO_SIGNED(478,11),
TO_SIGNED(441,11),
TO_SIGNED(402,11),
TO_SIGNED(362,11),
TO_SIGNED(320,11),
TO_SIGNED(276,11),
TO_SIGNED(232,11),
TO_SIGNED(187,11),
TO_SIGNED(141,11),
TO_SIGNED(95,11),
TO_SIGNED(48,11),
TO_SIGNED(1,11),
TO_SIGNED(-46,11),
TO_SIGNED(-93,11),
TO_SIGNED(-139,11),
TO_SIGNED(-185,11),
TO_SIGNED(-230,11),
TO_SIGNED(-275,11),
TO_SIGNED(-318,11),
TO_SIGNED(-360,11),
TO_SIGNED(-400,11),
TO_SIGNED(-439,11),
TO_SIGNED(-476,11),
TO_SIGNED(-512,11),
TO_SIGNED(-545,11),
TO_SIGNED(-576,11),
TO_SIGNED(-605,11),
TO_SIGNED(-632,11),
TO_SIGNED(-656,11),
TO_SIGNED(-677,11),
TO_SIGNED(-696,11),
TO_SIGNED(-712,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-715,11),
TO_SIGNED(-699,11),
TO_SIGNED(-681,11),
TO_SIGNED(-659,11),
TO_SIGNED(-636,11),
TO_SIGNED(-610,11),
TO_SIGNED(-581,11),
TO_SIGNED(-550,11),
TO_SIGNED(-517,11),
TO_SIGNED(-482,11),
TO_SIGNED(-445,11),
TO_SIGNED(-406,11),
TO_SIGNED(-366,11),
TO_SIGNED(-324,11),
TO_SIGNED(-281,11),
TO_SIGNED(-237,11),
TO_SIGNED(-192,11),
TO_SIGNED(-147,11),
TO_SIGNED(-100,11),
TO_SIGNED(-53,11),
TO_SIGNED(-6,11),
TO_SIGNED(41,11),
TO_SIGNED(87,11),
TO_SIGNED(134,11),
TO_SIGNED(180,11),
TO_SIGNED(225,11),
TO_SIGNED(270,11),
TO_SIGNED(313,11),
TO_SIGNED(355,11),
TO_SIGNED(396,11),
TO_SIGNED(435,11),
TO_SIGNED(472,11),
TO_SIGNED(508,11),
TO_SIGNED(541,11),
TO_SIGNED(573,11),
TO_SIGNED(602,11),
TO_SIGNED(629,11),
TO_SIGNED(653,11),
TO_SIGNED(675,11),
TO_SIGNED(694,11),
TO_SIGNED(711,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(729,11),
TO_SIGNED(716,11),
TO_SIGNED(701,11),
TO_SIGNED(683,11),
TO_SIGNED(662,11),
TO_SIGNED(639,11),
TO_SIGNED(613,11),
TO_SIGNED(584,11),
TO_SIGNED(554,11),
TO_SIGNED(521,11),
TO_SIGNED(486,11),
TO_SIGNED(449,11),
TO_SIGNED(411,11),
TO_SIGNED(371,11),
TO_SIGNED(329,11),
TO_SIGNED(286,11),
TO_SIGNED(242,11),
TO_SIGNED(197,11),
TO_SIGNED(152,11),
TO_SIGNED(105,11),
TO_SIGNED(59,11),
TO_SIGNED(12,11),
TO_SIGNED(-35,11),
TO_SIGNED(-82,11),
TO_SIGNED(-129,11),
TO_SIGNED(-175,11),
TO_SIGNED(-220,11),
TO_SIGNED(-265,11),
TO_SIGNED(-308,11),
TO_SIGNED(-350,11),
TO_SIGNED(-391,11),
TO_SIGNED(-430,11),
TO_SIGNED(-468,11),
TO_SIGNED(-504,11),
TO_SIGNED(-538,11),
TO_SIGNED(-569,11),
TO_SIGNED(-599,11),
TO_SIGNED(-626,11),
TO_SIGNED(-651,11),
TO_SIGNED(-673,11),
TO_SIGNED(-692,11),
TO_SIGNED(-709,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-685,11),
TO_SIGNED(-664,11),
TO_SIGNED(-641,11),
TO_SIGNED(-616,11),
TO_SIGNED(-588,11),
TO_SIGNED(-557,11),
TO_SIGNED(-525,11),
TO_SIGNED(-490,11),
TO_SIGNED(-454,11),
TO_SIGNED(-415,11),
TO_SIGNED(-375,11),
TO_SIGNED(-334,11),
TO_SIGNED(-291,11),
TO_SIGNED(-247,11),
TO_SIGNED(-203,11),
TO_SIGNED(-157,11),
TO_SIGNED(-111,11),
TO_SIGNED(-64,11),
TO_SIGNED(-17,11),
TO_SIGNED(30,11),
TO_SIGNED(77,11),
TO_SIGNED(123,11),
TO_SIGNED(169,11),
TO_SIGNED(215,11),
TO_SIGNED(260,11),
TO_SIGNED(303,11),
TO_SIGNED(345,11),
TO_SIGNED(387,11),
TO_SIGNED(426,11),
TO_SIGNED(464,11),
TO_SIGNED(500,11),
TO_SIGNED(534,11),
TO_SIGNED(566,11),
TO_SIGNED(596,11),
TO_SIGNED(623,11),
TO_SIGNED(648,11),
TO_SIGNED(670,11),
TO_SIGNED(690,11),
TO_SIGNED(707,11),
TO_SIGNED(721,11),
TO_SIGNED(733,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(705,11),
TO_SIGNED(687,11),
TO_SIGNED(667,11),
TO_SIGNED(644,11),
TO_SIGNED(619,11),
TO_SIGNED(591,11),
TO_SIGNED(561,11),
TO_SIGNED(529,11),
TO_SIGNED(494,11),
TO_SIGNED(458,11),
TO_SIGNED(420,11),
TO_SIGNED(380,11),
TO_SIGNED(339,11),
TO_SIGNED(296,11),
TO_SIGNED(252,11),
TO_SIGNED(208,11),
TO_SIGNED(162,11),
TO_SIGNED(116,11),
TO_SIGNED(69,11),
TO_SIGNED(22,11),
TO_SIGNED(-25,11),
TO_SIGNED(-71,11),
TO_SIGNED(-118,11),
TO_SIGNED(-164,11),
TO_SIGNED(-210,11),
TO_SIGNED(-255,11),
TO_SIGNED(-298,11),
TO_SIGNED(-341,11),
TO_SIGNED(-382,11),
TO_SIGNED(-422,11),
TO_SIGNED(-460,11),
TO_SIGNED(-496,11),
TO_SIGNED(-530,11),
TO_SIGNED(-562,11),
TO_SIGNED(-592,11),
TO_SIGNED(-620,11),
TO_SIGNED(-645,11),
TO_SIGNED(-668,11),
TO_SIGNED(-688,11),
TO_SIGNED(-705,11),
TO_SIGNED(-720,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-721,11),
TO_SIGNED(-706,11),
TO_SIGNED(-689,11),
TO_SIGNED(-669,11),
TO_SIGNED(-647,11),
TO_SIGNED(-622,11),
TO_SIGNED(-594,11),
TO_SIGNED(-564,11),
TO_SIGNED(-532,11),
TO_SIGNED(-498,11),
TO_SIGNED(-462,11),
TO_SIGNED(-424,11),
TO_SIGNED(-385,11),
TO_SIGNED(-344,11),
TO_SIGNED(-301,11),
TO_SIGNED(-258,11),
TO_SIGNED(-213,11),
TO_SIGNED(-167,11),
TO_SIGNED(-121,11),
TO_SIGNED(-75,11),
TO_SIGNED(-28,11),
TO_SIGNED(19,11),
TO_SIGNED(66,11),
TO_SIGNED(113,11),
TO_SIGNED(159,11),
TO_SIGNED(205,11),
TO_SIGNED(249,11),
TO_SIGNED(293,11),
TO_SIGNED(336,11),
TO_SIGNED(377,11),
TO_SIGNED(417,11),
TO_SIGNED(455,11),
TO_SIGNED(492,11),
TO_SIGNED(526,11),
TO_SIGNED(559,11),
TO_SIGNED(589,11),
TO_SIGNED(617,11),
TO_SIGNED(642,11),
TO_SIGNED(665,11),
TO_SIGNED(686,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(708,11),
TO_SIGNED(691,11),
TO_SIGNED(672,11),
TO_SIGNED(650,11),
TO_SIGNED(625,11),
TO_SIGNED(598,11),
TO_SIGNED(568,11),
TO_SIGNED(536,11),
TO_SIGNED(502,11),
TO_SIGNED(466,11),
TO_SIGNED(429,11),
TO_SIGNED(389,11),
TO_SIGNED(348,11),
TO_SIGNED(306,11),
TO_SIGNED(263,11),
TO_SIGNED(218,11),
TO_SIGNED(173,11),
TO_SIGNED(127,11),
TO_SIGNED(80,11),
TO_SIGNED(33,11),
TO_SIGNED(-14,11),
TO_SIGNED(-61,11),
TO_SIGNED(-108,11),
TO_SIGNED(-154,11),
TO_SIGNED(-200,11),
TO_SIGNED(-244,11),
TO_SIGNED(-288,11),
TO_SIGNED(-331,11),
TO_SIGNED(-373,11),
TO_SIGNED(-413,11),
TO_SIGNED(-451,11),
TO_SIGNED(-488,11),
TO_SIGNED(-523,11),
TO_SIGNED(-555,11),
TO_SIGNED(-586,11),
TO_SIGNED(-614,11),
TO_SIGNED(-640,11),
TO_SIGNED(-663,11),
TO_SIGNED(-684,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-729,11),
TO_SIGNED(-739,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-710,11),
TO_SIGNED(-693,11),
TO_SIGNED(-674,11),
TO_SIGNED(-652,11),
TO_SIGNED(-628,11),
TO_SIGNED(-601,11),
TO_SIGNED(-571,11),
TO_SIGNED(-540,11),
TO_SIGNED(-506,11),
TO_SIGNED(-471,11),
TO_SIGNED(-433,11),
TO_SIGNED(-394,11),
TO_SIGNED(-353,11),
TO_SIGNED(-311,11),
TO_SIGNED(-268,11),
TO_SIGNED(-223,11),
TO_SIGNED(-178,11),
TO_SIGNED(-132,11),
TO_SIGNED(-85,11),
TO_SIGNED(-38,11),
TO_SIGNED(9,11),
TO_SIGNED(56,11),
TO_SIGNED(102,11),
TO_SIGNED(149,11),
TO_SIGNED(194,11),
TO_SIGNED(239,11),
TO_SIGNED(283,11),
TO_SIGNED(326,11),
TO_SIGNED(368,11),
TO_SIGNED(408,11),
TO_SIGNED(447,11),
TO_SIGNED(484,11),
TO_SIGNED(519,11),
TO_SIGNED(552,11),
TO_SIGNED(582,11),
TO_SIGNED(611,11),
TO_SIGNED(637,11),
TO_SIGNED(660,11),
TO_SIGNED(681,11),
TO_SIGNED(700,11),
TO_SIGNED(715,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(736,11),
TO_SIGNED(725,11),
TO_SIGNED(712,11),
TO_SIGNED(695,11),
TO_SIGNED(676,11),
TO_SIGNED(655,11),
TO_SIGNED(631,11),
TO_SIGNED(604,11),
TO_SIGNED(575,11),
TO_SIGNED(544,11),
TO_SIGNED(510,11),
TO_SIGNED(475,11),
TO_SIGNED(437,11),
TO_SIGNED(398,11),
TO_SIGNED(358,11),
TO_SIGNED(316,11),
TO_SIGNED(273,11),
TO_SIGNED(228,11),
TO_SIGNED(183,11),
TO_SIGNED(137,11),
TO_SIGNED(91,11),
TO_SIGNED(44,11),
TO_SIGNED(-3,11),
TO_SIGNED(-50,11),
TO_SIGNED(-97,11),
TO_SIGNED(-143,11),
TO_SIGNED(-189,11),
TO_SIGNED(-234,11),
TO_SIGNED(-278,11),
TO_SIGNED(-322,11),
TO_SIGNED(-363,11),
TO_SIGNED(-404,11),
TO_SIGNED(-443,11),
TO_SIGNED(-480,11),
TO_SIGNED(-515,11),
TO_SIGNED(-548,11),
TO_SIGNED(-579,11),
TO_SIGNED(-608,11),
TO_SIGNED(-634,11),
TO_SIGNED(-658,11),
TO_SIGNED(-679,11),
TO_SIGNED(-698,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-679,11),
TO_SIGNED(-657,11),
TO_SIGNED(-633,11),
TO_SIGNED(-607,11),
TO_SIGNED(-578,11),
TO_SIGNED(-547,11),
TO_SIGNED(-514,11),
TO_SIGNED(-479,11),
TO_SIGNED(-442,11),
TO_SIGNED(-403,11),
TO_SIGNED(-362,11),
TO_SIGNED(-321,11),
TO_SIGNED(-277,11),
TO_SIGNED(-233,11),
TO_SIGNED(-188,11),
TO_SIGNED(-142,11),
TO_SIGNED(-96,11),
TO_SIGNED(-49,11),
TO_SIGNED(-2,11),
TO_SIGNED(45,11),
TO_SIGNED(92,11),
TO_SIGNED(138,11),
TO_SIGNED(184,11),
TO_SIGNED(229,11),
TO_SIGNED(274,11),
TO_SIGNED(317,11),
TO_SIGNED(359,11),
TO_SIGNED(399,11),
TO_SIGNED(438,11),
TO_SIGNED(476,11),
TO_SIGNED(511,11),
TO_SIGNED(544,11),
TO_SIGNED(576,11),
TO_SIGNED(605,11),
TO_SIGNED(631,11),
TO_SIGNED(655,11),
TO_SIGNED(677,11),
TO_SIGNED(696,11),
TO_SIGNED(712,11),
TO_SIGNED(725,11),
TO_SIGNED(736,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(715,11),
TO_SIGNED(699,11),
TO_SIGNED(681,11),
TO_SIGNED(660,11),
TO_SIGNED(636,11),
TO_SIGNED(610,11),
TO_SIGNED(582,11),
TO_SIGNED(551,11),
TO_SIGNED(518,11),
TO_SIGNED(483,11),
TO_SIGNED(446,11),
TO_SIGNED(407,11),
TO_SIGNED(367,11),
TO_SIGNED(325,11),
TO_SIGNED(282,11),
TO_SIGNED(238,11),
TO_SIGNED(193,11),
TO_SIGNED(148,11),
TO_SIGNED(101,11),
TO_SIGNED(54,11),
TO_SIGNED(7,11),
TO_SIGNED(-40,11),
TO_SIGNED(-86,11),
TO_SIGNED(-133,11),
TO_SIGNED(-179,11),
TO_SIGNED(-224,11),
TO_SIGNED(-269,11),
TO_SIGNED(-312,11),
TO_SIGNED(-354,11),
TO_SIGNED(-395,11),
TO_SIGNED(-434,11),
TO_SIGNED(-471,11),
TO_SIGNED(-507,11),
TO_SIGNED(-541,11),
TO_SIGNED(-572,11),
TO_SIGNED(-601,11),
TO_SIGNED(-628,11),
TO_SIGNED(-653,11),
TO_SIGNED(-675,11),
TO_SIGNED(-694,11),
TO_SIGNED(-710,11),
TO_SIGNED(-724,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-701,11),
TO_SIGNED(-683,11),
TO_SIGNED(-662,11),
TO_SIGNED(-639,11),
TO_SIGNED(-613,11),
TO_SIGNED(-585,11),
TO_SIGNED(-554,11),
TO_SIGNED(-522,11),
TO_SIGNED(-487,11),
TO_SIGNED(-450,11),
TO_SIGNED(-412,11),
TO_SIGNED(-372,11),
TO_SIGNED(-330,11),
TO_SIGNED(-287,11),
TO_SIGNED(-243,11),
TO_SIGNED(-198,11),
TO_SIGNED(-153,11),
TO_SIGNED(-106,11),
TO_SIGNED(-60,11),
TO_SIGNED(-13,11),
TO_SIGNED(34,11),
TO_SIGNED(81,11),
TO_SIGNED(128,11),
TO_SIGNED(174,11),
TO_SIGNED(219,11),
TO_SIGNED(264,11),
TO_SIGNED(307,11),
TO_SIGNED(349,11),
TO_SIGNED(390,11),
TO_SIGNED(430,11),
TO_SIGNED(467,11),
TO_SIGNED(503,11),
TO_SIGNED(537,11),
TO_SIGNED(569,11),
TO_SIGNED(598,11),
TO_SIGNED(625,11),
TO_SIGNED(650,11),
TO_SIGNED(672,11),
TO_SIGNED(692,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(730,11),
TO_SIGNED(718,11),
TO_SIGNED(703,11),
TO_SIGNED(685,11),
TO_SIGNED(665,11),
TO_SIGNED(642,11),
TO_SIGNED(616,11),
TO_SIGNED(588,11),
TO_SIGNED(558,11),
TO_SIGNED(526,11),
TO_SIGNED(491,11),
TO_SIGNED(455,11),
TO_SIGNED(416,11),
TO_SIGNED(376,11),
TO_SIGNED(335,11),
TO_SIGNED(292,11),
TO_SIGNED(248,11),
TO_SIGNED(204,11),
TO_SIGNED(158,11),
TO_SIGNED(112,11),
TO_SIGNED(65,11),
TO_SIGNED(18,11),
TO_SIGNED(-29,11),
TO_SIGNED(-76,11),
TO_SIGNED(-122,11),
TO_SIGNED(-168,11),
TO_SIGNED(-214,11),
TO_SIGNED(-259,11),
TO_SIGNED(-302,11),
TO_SIGNED(-345,11),
TO_SIGNED(-386,11),
TO_SIGNED(-425,11),
TO_SIGNED(-463,11),
TO_SIGNED(-499,11),
TO_SIGNED(-533,11),
TO_SIGNED(-565,11),
TO_SIGNED(-595,11),
TO_SIGNED(-622,11),
TO_SIGNED(-647,11),
TO_SIGNED(-670,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-721,11),
TO_SIGNED(-733,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-720,11),
TO_SIGNED(-705,11),
TO_SIGNED(-688,11),
TO_SIGNED(-667,11),
TO_SIGNED(-645,11),
TO_SIGNED(-619,11),
TO_SIGNED(-592,11),
TO_SIGNED(-562,11),
TO_SIGNED(-529,11),
TO_SIGNED(-495,11),
TO_SIGNED(-459,11),
TO_SIGNED(-421,11),
TO_SIGNED(-381,11),
TO_SIGNED(-340,11),
TO_SIGNED(-297,11),
TO_SIGNED(-254,11),
TO_SIGNED(-209,11),
TO_SIGNED(-163,11),
TO_SIGNED(-117,11),
TO_SIGNED(-70,11),
TO_SIGNED(-24,11),
TO_SIGNED(24,11),
TO_SIGNED(70,11),
TO_SIGNED(117,11),
TO_SIGNED(163,11),
TO_SIGNED(209,11),
TO_SIGNED(254,11),
TO_SIGNED(297,11),
TO_SIGNED(340,11),
TO_SIGNED(381,11),
TO_SIGNED(421,11),
TO_SIGNED(459,11),
TO_SIGNED(495,11),
TO_SIGNED(529,11),
TO_SIGNED(562,11),
TO_SIGNED(592,11),
TO_SIGNED(619,11),
TO_SIGNED(645,11),
TO_SIGNED(667,11),
TO_SIGNED(688,11),
TO_SIGNED(705,11),
TO_SIGNED(720,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(733,11),
TO_SIGNED(721,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(670,11),
TO_SIGNED(647,11),
TO_SIGNED(622,11),
TO_SIGNED(595,11),
TO_SIGNED(565,11),
TO_SIGNED(533,11),
TO_SIGNED(499,11),
TO_SIGNED(463,11),
TO_SIGNED(425,11),
TO_SIGNED(386,11),
TO_SIGNED(345,11),
TO_SIGNED(302,11),
TO_SIGNED(259,11),
TO_SIGNED(214,11),
TO_SIGNED(168,11),
TO_SIGNED(122,11),
TO_SIGNED(76,11),
TO_SIGNED(29,11),
TO_SIGNED(-18,11),
TO_SIGNED(-65,11),
TO_SIGNED(-112,11),
TO_SIGNED(-158,11),
TO_SIGNED(-204,11),
TO_SIGNED(-248,11),
TO_SIGNED(-292,11),
TO_SIGNED(-335,11),
TO_SIGNED(-376,11),
TO_SIGNED(-416,11),
TO_SIGNED(-455,11),
TO_SIGNED(-491,11),
TO_SIGNED(-526,11),
TO_SIGNED(-558,11),
TO_SIGNED(-588,11),
TO_SIGNED(-616,11),
TO_SIGNED(-642,11),
TO_SIGNED(-665,11),
TO_SIGNED(-685,11),
TO_SIGNED(-703,11),
TO_SIGNED(-718,11),
TO_SIGNED(-730,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-692,11),
TO_SIGNED(-672,11),
TO_SIGNED(-650,11),
TO_SIGNED(-625,11),
TO_SIGNED(-598,11),
TO_SIGNED(-569,11),
TO_SIGNED(-537,11),
TO_SIGNED(-503,11),
TO_SIGNED(-467,11),
TO_SIGNED(-430,11),
TO_SIGNED(-390,11),
TO_SIGNED(-349,11),
TO_SIGNED(-307,11),
TO_SIGNED(-264,11),
TO_SIGNED(-219,11),
TO_SIGNED(-174,11),
TO_SIGNED(-128,11),
TO_SIGNED(-81,11),
TO_SIGNED(-34,11),
TO_SIGNED(13,11),
TO_SIGNED(60,11),
TO_SIGNED(106,11),
TO_SIGNED(153,11),
TO_SIGNED(198,11),
TO_SIGNED(243,11),
TO_SIGNED(287,11),
TO_SIGNED(330,11),
TO_SIGNED(372,11),
TO_SIGNED(412,11),
TO_SIGNED(450,11),
TO_SIGNED(487,11),
TO_SIGNED(522,11),
TO_SIGNED(554,11),
TO_SIGNED(585,11),
TO_SIGNED(613,11),
TO_SIGNED(639,11),
TO_SIGNED(662,11),
TO_SIGNED(683,11),
TO_SIGNED(701,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(724,11),
TO_SIGNED(710,11),
TO_SIGNED(694,11),
TO_SIGNED(675,11),
TO_SIGNED(653,11),
TO_SIGNED(628,11),
TO_SIGNED(601,11),
TO_SIGNED(572,11),
TO_SIGNED(541,11),
TO_SIGNED(507,11),
TO_SIGNED(471,11),
TO_SIGNED(434,11),
TO_SIGNED(395,11),
TO_SIGNED(354,11),
TO_SIGNED(312,11),
TO_SIGNED(269,11),
TO_SIGNED(224,11),
TO_SIGNED(179,11),
TO_SIGNED(133,11),
TO_SIGNED(86,11),
TO_SIGNED(40,11),
TO_SIGNED(-7,11),
TO_SIGNED(-54,11),
TO_SIGNED(-101,11),
TO_SIGNED(-148,11),
TO_SIGNED(-193,11),
TO_SIGNED(-238,11),
TO_SIGNED(-282,11),
TO_SIGNED(-325,11),
TO_SIGNED(-367,11),
TO_SIGNED(-407,11),
TO_SIGNED(-446,11),
TO_SIGNED(-483,11),
TO_SIGNED(-518,11),
TO_SIGNED(-551,11),
TO_SIGNED(-582,11),
TO_SIGNED(-610,11),
TO_SIGNED(-636,11),
TO_SIGNED(-660,11),
TO_SIGNED(-681,11),
TO_SIGNED(-699,11),
TO_SIGNED(-715,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-736,11),
TO_SIGNED(-725,11),
TO_SIGNED(-712,11),
TO_SIGNED(-696,11),
TO_SIGNED(-677,11),
TO_SIGNED(-655,11),
TO_SIGNED(-631,11),
TO_SIGNED(-605,11),
TO_SIGNED(-576,11),
TO_SIGNED(-544,11),
TO_SIGNED(-511,11),
TO_SIGNED(-476,11),
TO_SIGNED(-438,11),
TO_SIGNED(-399,11),
TO_SIGNED(-359,11),
TO_SIGNED(-317,11),
TO_SIGNED(-274,11),
TO_SIGNED(-229,11),
TO_SIGNED(-184,11),
TO_SIGNED(-138,11),
TO_SIGNED(-92,11),
TO_SIGNED(-45,11),
TO_SIGNED(2,11),
TO_SIGNED(49,11),
TO_SIGNED(96,11),
TO_SIGNED(142,11),
TO_SIGNED(188,11),
TO_SIGNED(233,11),
TO_SIGNED(277,11),
TO_SIGNED(321,11),
TO_SIGNED(362,11),
TO_SIGNED(403,11),
TO_SIGNED(442,11),
TO_SIGNED(479,11),
TO_SIGNED(514,11),
TO_SIGNED(547,11),
TO_SIGNED(578,11),
TO_SIGNED(607,11),
TO_SIGNED(633,11),
TO_SIGNED(657,11),
TO_SIGNED(679,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(698,11),
TO_SIGNED(679,11),
TO_SIGNED(658,11),
TO_SIGNED(634,11),
TO_SIGNED(608,11),
TO_SIGNED(579,11),
TO_SIGNED(548,11),
TO_SIGNED(515,11),
TO_SIGNED(480,11),
TO_SIGNED(443,11),
TO_SIGNED(404,11),
TO_SIGNED(363,11),
TO_SIGNED(322,11),
TO_SIGNED(278,11),
TO_SIGNED(234,11),
TO_SIGNED(189,11),
TO_SIGNED(143,11),
TO_SIGNED(97,11),
TO_SIGNED(50,11),
TO_SIGNED(3,11),
TO_SIGNED(-44,11),
TO_SIGNED(-91,11),
TO_SIGNED(-137,11),
TO_SIGNED(-183,11),
TO_SIGNED(-228,11),
TO_SIGNED(-273,11),
TO_SIGNED(-316,11),
TO_SIGNED(-358,11),
TO_SIGNED(-398,11),
TO_SIGNED(-437,11),
TO_SIGNED(-475,11),
TO_SIGNED(-510,11),
TO_SIGNED(-544,11),
TO_SIGNED(-575,11),
TO_SIGNED(-604,11),
TO_SIGNED(-631,11),
TO_SIGNED(-655,11),
TO_SIGNED(-676,11),
TO_SIGNED(-695,11),
TO_SIGNED(-712,11),
TO_SIGNED(-725,11),
TO_SIGNED(-736,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-715,11),
TO_SIGNED(-700,11),
TO_SIGNED(-681,11),
TO_SIGNED(-660,11),
TO_SIGNED(-637,11),
TO_SIGNED(-611,11),
TO_SIGNED(-582,11),
TO_SIGNED(-552,11),
TO_SIGNED(-519,11),
TO_SIGNED(-484,11),
TO_SIGNED(-447,11),
TO_SIGNED(-408,11),
TO_SIGNED(-368,11),
TO_SIGNED(-326,11),
TO_SIGNED(-283,11),
TO_SIGNED(-239,11),
TO_SIGNED(-194,11),
TO_SIGNED(-149,11),
TO_SIGNED(-102,11),
TO_SIGNED(-56,11),
TO_SIGNED(-9,11),
TO_SIGNED(38,11),
TO_SIGNED(85,11),
TO_SIGNED(132,11),
TO_SIGNED(178,11),
TO_SIGNED(223,11),
TO_SIGNED(268,11),
TO_SIGNED(311,11),
TO_SIGNED(353,11),
TO_SIGNED(394,11),
TO_SIGNED(433,11),
TO_SIGNED(471,11),
TO_SIGNED(506,11),
TO_SIGNED(540,11),
TO_SIGNED(571,11),
TO_SIGNED(601,11),
TO_SIGNED(628,11),
TO_SIGNED(652,11),
TO_SIGNED(674,11),
TO_SIGNED(693,11),
TO_SIGNED(710,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(739,11),
TO_SIGNED(729,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(684,11),
TO_SIGNED(663,11),
TO_SIGNED(640,11),
TO_SIGNED(614,11),
TO_SIGNED(586,11),
TO_SIGNED(555,11),
TO_SIGNED(523,11),
TO_SIGNED(488,11),
TO_SIGNED(451,11),
TO_SIGNED(413,11),
TO_SIGNED(373,11),
TO_SIGNED(331,11),
TO_SIGNED(288,11),
TO_SIGNED(244,11),
TO_SIGNED(200,11),
TO_SIGNED(154,11),
TO_SIGNED(108,11),
TO_SIGNED(61,11),
TO_SIGNED(14,11),
TO_SIGNED(-33,11),
TO_SIGNED(-80,11),
TO_SIGNED(-127,11),
TO_SIGNED(-173,11),
TO_SIGNED(-218,11),
TO_SIGNED(-263,11),
TO_SIGNED(-306,11),
TO_SIGNED(-348,11),
TO_SIGNED(-389,11),
TO_SIGNED(-429,11),
TO_SIGNED(-466,11),
TO_SIGNED(-502,11),
TO_SIGNED(-536,11),
TO_SIGNED(-568,11),
TO_SIGNED(-598,11),
TO_SIGNED(-625,11),
TO_SIGNED(-650,11),
TO_SIGNED(-672,11),
TO_SIGNED(-691,11),
TO_SIGNED(-708,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-686,11),
TO_SIGNED(-665,11),
TO_SIGNED(-642,11),
TO_SIGNED(-617,11),
TO_SIGNED(-589,11),
TO_SIGNED(-559,11),
TO_SIGNED(-526,11),
TO_SIGNED(-492,11),
TO_SIGNED(-455,11),
TO_SIGNED(-417,11),
TO_SIGNED(-377,11),
TO_SIGNED(-336,11),
TO_SIGNED(-293,11),
TO_SIGNED(-249,11),
TO_SIGNED(-205,11),
TO_SIGNED(-159,11),
TO_SIGNED(-113,11),
TO_SIGNED(-66,11),
TO_SIGNED(-19,11),
TO_SIGNED(28,11),
TO_SIGNED(75,11),
TO_SIGNED(121,11),
TO_SIGNED(167,11),
TO_SIGNED(213,11),
TO_SIGNED(258,11),
TO_SIGNED(301,11),
TO_SIGNED(344,11),
TO_SIGNED(385,11),
TO_SIGNED(424,11),
TO_SIGNED(462,11),
TO_SIGNED(498,11),
TO_SIGNED(532,11),
TO_SIGNED(564,11),
TO_SIGNED(594,11),
TO_SIGNED(622,11),
TO_SIGNED(647,11),
TO_SIGNED(669,11),
TO_SIGNED(689,11),
TO_SIGNED(706,11),
TO_SIGNED(721,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(720,11),
TO_SIGNED(705,11),
TO_SIGNED(688,11),
TO_SIGNED(668,11),
TO_SIGNED(645,11),
TO_SIGNED(620,11),
TO_SIGNED(592,11),
TO_SIGNED(562,11),
TO_SIGNED(530,11),
TO_SIGNED(496,11),
TO_SIGNED(460,11),
TO_SIGNED(422,11),
TO_SIGNED(382,11),
TO_SIGNED(341,11),
TO_SIGNED(298,11),
TO_SIGNED(255,11),
TO_SIGNED(210,11),
TO_SIGNED(164,11),
TO_SIGNED(118,11),
TO_SIGNED(71,11),
TO_SIGNED(25,11),
TO_SIGNED(-22,11),
TO_SIGNED(-69,11),
TO_SIGNED(-116,11),
TO_SIGNED(-162,11),
TO_SIGNED(-208,11),
TO_SIGNED(-252,11),
TO_SIGNED(-296,11),
TO_SIGNED(-339,11),
TO_SIGNED(-380,11),
TO_SIGNED(-420,11),
TO_SIGNED(-458,11),
TO_SIGNED(-494,11),
TO_SIGNED(-529,11),
TO_SIGNED(-561,11),
TO_SIGNED(-591,11),
TO_SIGNED(-619,11),
TO_SIGNED(-644,11),
TO_SIGNED(-667,11),
TO_SIGNED(-687,11),
TO_SIGNED(-705,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-733,11),
TO_SIGNED(-721,11),
TO_SIGNED(-707,11),
TO_SIGNED(-690,11),
TO_SIGNED(-670,11),
TO_SIGNED(-648,11),
TO_SIGNED(-623,11),
TO_SIGNED(-596,11),
TO_SIGNED(-566,11),
TO_SIGNED(-534,11),
TO_SIGNED(-500,11),
TO_SIGNED(-464,11),
TO_SIGNED(-426,11),
TO_SIGNED(-387,11),
TO_SIGNED(-345,11),
TO_SIGNED(-303,11),
TO_SIGNED(-260,11),
TO_SIGNED(-215,11),
TO_SIGNED(-169,11),
TO_SIGNED(-123,11),
TO_SIGNED(-77,11),
TO_SIGNED(-30,11),
TO_SIGNED(17,11),
TO_SIGNED(64,11),
TO_SIGNED(111,11),
TO_SIGNED(157,11),
TO_SIGNED(203,11),
TO_SIGNED(247,11),
TO_SIGNED(291,11),
TO_SIGNED(334,11),
TO_SIGNED(375,11),
TO_SIGNED(415,11),
TO_SIGNED(454,11),
TO_SIGNED(490,11),
TO_SIGNED(525,11),
TO_SIGNED(557,11),
TO_SIGNED(588,11),
TO_SIGNED(616,11),
TO_SIGNED(641,11),
TO_SIGNED(664,11),
TO_SIGNED(685,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(709,11),
TO_SIGNED(692,11),
TO_SIGNED(673,11),
TO_SIGNED(651,11),
TO_SIGNED(626,11),
TO_SIGNED(599,11),
TO_SIGNED(569,11),
TO_SIGNED(538,11),
TO_SIGNED(504,11),
TO_SIGNED(468,11),
TO_SIGNED(430,11),
TO_SIGNED(391,11),
TO_SIGNED(350,11),
TO_SIGNED(308,11),
TO_SIGNED(265,11),
TO_SIGNED(220,11),
TO_SIGNED(175,11),
TO_SIGNED(129,11),
TO_SIGNED(82,11),
TO_SIGNED(35,11),
TO_SIGNED(-12,11),
TO_SIGNED(-59,11),
TO_SIGNED(-105,11),
TO_SIGNED(-152,11),
TO_SIGNED(-197,11),
TO_SIGNED(-242,11),
TO_SIGNED(-286,11),
TO_SIGNED(-329,11),
TO_SIGNED(-371,11),
TO_SIGNED(-411,11),
TO_SIGNED(-449,11),
TO_SIGNED(-486,11),
TO_SIGNED(-521,11),
TO_SIGNED(-554,11),
TO_SIGNED(-584,11),
TO_SIGNED(-613,11),
TO_SIGNED(-639,11),
TO_SIGNED(-662,11),
TO_SIGNED(-683,11),
TO_SIGNED(-701,11),
TO_SIGNED(-716,11),
TO_SIGNED(-729,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-711,11),
TO_SIGNED(-694,11),
TO_SIGNED(-675,11),
TO_SIGNED(-653,11),
TO_SIGNED(-629,11),
TO_SIGNED(-602,11),
TO_SIGNED(-573,11),
TO_SIGNED(-541,11),
TO_SIGNED(-508,11),
TO_SIGNED(-472,11),
TO_SIGNED(-435,11),
TO_SIGNED(-396,11),
TO_SIGNED(-355,11),
TO_SIGNED(-313,11),
TO_SIGNED(-270,11),
TO_SIGNED(-225,11),
TO_SIGNED(-180,11),
TO_SIGNED(-134,11),
TO_SIGNED(-87,11),
TO_SIGNED(-41,11),
TO_SIGNED(6,11),
TO_SIGNED(53,11),
TO_SIGNED(100,11),
TO_SIGNED(147,11),
TO_SIGNED(192,11),
TO_SIGNED(237,11),
TO_SIGNED(281,11),
TO_SIGNED(324,11),
TO_SIGNED(366,11),
TO_SIGNED(406,11),
TO_SIGNED(445,11),
TO_SIGNED(482,11),
TO_SIGNED(517,11),
TO_SIGNED(550,11),
TO_SIGNED(581,11),
TO_SIGNED(610,11),
TO_SIGNED(636,11),
TO_SIGNED(659,11),
TO_SIGNED(681,11),
TO_SIGNED(699,11),
TO_SIGNED(715,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(712,11),
TO_SIGNED(696,11),
TO_SIGNED(677,11),
TO_SIGNED(656,11),
TO_SIGNED(632,11),
TO_SIGNED(605,11),
TO_SIGNED(576,11),
TO_SIGNED(545,11),
TO_SIGNED(512,11),
TO_SIGNED(476,11),
TO_SIGNED(439,11),
TO_SIGNED(400,11),
TO_SIGNED(360,11),
TO_SIGNED(318,11),
TO_SIGNED(275,11),
TO_SIGNED(230,11),
TO_SIGNED(185,11),
TO_SIGNED(139,11),
TO_SIGNED(93,11),
TO_SIGNED(46,11),
TO_SIGNED(-1,11),
TO_SIGNED(-48,11),
TO_SIGNED(-95,11),
TO_SIGNED(-141,11),
TO_SIGNED(-187,11),
TO_SIGNED(-232,11),
TO_SIGNED(-276,11),
TO_SIGNED(-320,11),
TO_SIGNED(-362,11),
TO_SIGNED(-402,11),
TO_SIGNED(-441,11),
TO_SIGNED(-478,11),
TO_SIGNED(-513,11),
TO_SIGNED(-547,11),
TO_SIGNED(-578,11),
TO_SIGNED(-606,11),
TO_SIGNED(-633,11),
TO_SIGNED(-657,11),
TO_SIGNED(-678,11),
TO_SIGNED(-697,11),
TO_SIGNED(-713,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-714,11),
TO_SIGNED(-698,11),
TO_SIGNED(-680,11),
TO_SIGNED(-658,11),
TO_SIGNED(-635,11),
TO_SIGNED(-608,11),
TO_SIGNED(-580,11),
TO_SIGNED(-549,11),
TO_SIGNED(-516,11),
TO_SIGNED(-480,11),
TO_SIGNED(-443,11),
TO_SIGNED(-405,11),
TO_SIGNED(-364,11),
TO_SIGNED(-323,11),
TO_SIGNED(-279,11),
TO_SIGNED(-235,11),
TO_SIGNED(-190,11),
TO_SIGNED(-144,11),
TO_SIGNED(-98,11),
TO_SIGNED(-51,11),
TO_SIGNED(-4,11),
TO_SIGNED(43,11),
TO_SIGNED(90,11),
TO_SIGNED(136,11),
TO_SIGNED(182,11),
TO_SIGNED(227,11),
TO_SIGNED(272,11),
TO_SIGNED(315,11),
TO_SIGNED(357,11),
TO_SIGNED(397,11),
TO_SIGNED(437,11),
TO_SIGNED(474,11),
TO_SIGNED(509,11),
TO_SIGNED(543,11),
TO_SIGNED(574,11),
TO_SIGNED(603,11),
TO_SIGNED(630,11),
TO_SIGNED(654,11),
TO_SIGNED(676,11),
TO_SIGNED(695,11),
TO_SIGNED(711,11),
TO_SIGNED(725,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(716,11),
TO_SIGNED(700,11),
TO_SIGNED(682,11),
TO_SIGNED(661,11),
TO_SIGNED(637,11),
TO_SIGNED(611,11),
TO_SIGNED(583,11),
TO_SIGNED(552,11),
TO_SIGNED(519,11),
TO_SIGNED(485,11),
TO_SIGNED(448,11),
TO_SIGNED(409,11),
TO_SIGNED(369,11),
TO_SIGNED(327,11),
TO_SIGNED(284,11),
TO_SIGNED(240,11),
TO_SIGNED(195,11),
TO_SIGNED(150,11),
TO_SIGNED(103,11),
TO_SIGNED(57,11),
TO_SIGNED(10,11),
TO_SIGNED(-37,11),
TO_SIGNED(-84,11),
TO_SIGNED(-131,11),
TO_SIGNED(-177,11),
TO_SIGNED(-222,11),
TO_SIGNED(-267,11),
TO_SIGNED(-310,11),
TO_SIGNED(-352,11),
TO_SIGNED(-393,11),
TO_SIGNED(-432,11),
TO_SIGNED(-470,11),
TO_SIGNED(-505,11),
TO_SIGNED(-539,11),
TO_SIGNED(-571,11),
TO_SIGNED(-600,11),
TO_SIGNED(-627,11),
TO_SIGNED(-652,11),
TO_SIGNED(-674,11),
TO_SIGNED(-693,11),
TO_SIGNED(-710,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-702,11),
TO_SIGNED(-684,11),
TO_SIGNED(-663,11),
TO_SIGNED(-640,11),
TO_SIGNED(-615,11),
TO_SIGNED(-586,11),
TO_SIGNED(-556,11),
TO_SIGNED(-523,11),
TO_SIGNED(-489,11),
TO_SIGNED(-452,11),
TO_SIGNED(-414,11),
TO_SIGNED(-374,11),
TO_SIGNED(-332,11),
TO_SIGNED(-289,11),
TO_SIGNED(-245,11),
TO_SIGNED(-201,11),
TO_SIGNED(-155,11),
TO_SIGNED(-109,11),
TO_SIGNED(-62,11),
TO_SIGNED(-15,11),
TO_SIGNED(32,11),
TO_SIGNED(79,11),
TO_SIGNED(125,11),
TO_SIGNED(172,11),
TO_SIGNED(217,11),
TO_SIGNED(262,11),
TO_SIGNED(305,11),
TO_SIGNED(347,11),
TO_SIGNED(388,11),
TO_SIGNED(428,11),
TO_SIGNED(466,11),
TO_SIGNED(501,11),
TO_SIGNED(535,11),
TO_SIGNED(567,11),
TO_SIGNED(597,11),
TO_SIGNED(624,11),
TO_SIGNED(649,11),
TO_SIGNED(671,11),
TO_SIGNED(691,11),
TO_SIGNED(708,11),
TO_SIGNED(722,11),
TO_SIGNED(733,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(704,11),
TO_SIGNED(686,11),
TO_SIGNED(666,11),
TO_SIGNED(643,11),
TO_SIGNED(618,11),
TO_SIGNED(590,11),
TO_SIGNED(559,11),
TO_SIGNED(527,11),
TO_SIGNED(493,11),
TO_SIGNED(456,11),
TO_SIGNED(418,11),
TO_SIGNED(378,11),
TO_SIGNED(337,11),
TO_SIGNED(294,11),
TO_SIGNED(250,11),
TO_SIGNED(206,11),
TO_SIGNED(160,11),
TO_SIGNED(114,11),
TO_SIGNED(67,11),
TO_SIGNED(20,11),
TO_SIGNED(-27,11),
TO_SIGNED(-74,11),
TO_SIGNED(-120,11),
TO_SIGNED(-166,11),
TO_SIGNED(-212,11),
TO_SIGNED(-257,11),
TO_SIGNED(-300,11),
TO_SIGNED(-343,11),
TO_SIGNED(-384,11),
TO_SIGNED(-423,11),
TO_SIGNED(-461,11),
TO_SIGNED(-497,11),
TO_SIGNED(-532,11),
TO_SIGNED(-564,11),
TO_SIGNED(-594,11),
TO_SIGNED(-621,11),
TO_SIGNED(-646,11),
TO_SIGNED(-669,11),
TO_SIGNED(-689,11),
TO_SIGNED(-706,11),
TO_SIGNED(-721,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-720,11),
TO_SIGNED(-706,11),
TO_SIGNED(-688,11),
TO_SIGNED(-668,11),
TO_SIGNED(-646,11),
TO_SIGNED(-621,11),
TO_SIGNED(-593,11),
TO_SIGNED(-563,11),
TO_SIGNED(-531,11),
TO_SIGNED(-497,11),
TO_SIGNED(-460,11),
TO_SIGNED(-422,11),
TO_SIGNED(-383,11),
TO_SIGNED(-342,11),
TO_SIGNED(-299,11),
TO_SIGNED(-256,11),
TO_SIGNED(-211,11),
TO_SIGNED(-165,11),
TO_SIGNED(-119,11),
TO_SIGNED(-73,11),
TO_SIGNED(-26,11),
TO_SIGNED(21,11),
TO_SIGNED(68,11),
TO_SIGNED(115,11),
TO_SIGNED(161,11),
TO_SIGNED(207,11),
TO_SIGNED(251,11),
TO_SIGNED(295,11),
TO_SIGNED(338,11),
TO_SIGNED(379,11),
TO_SIGNED(419,11),
TO_SIGNED(457,11),
TO_SIGNED(493,11),
TO_SIGNED(528,11),
TO_SIGNED(560,11),
TO_SIGNED(590,11),
TO_SIGNED(618,11),
TO_SIGNED(644,11),
TO_SIGNED(666,11),
TO_SIGNED(687,11),
TO_SIGNED(704,11),
TO_SIGNED(719,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(671,11),
TO_SIGNED(648,11),
TO_SIGNED(624,11),
TO_SIGNED(596,11),
TO_SIGNED(567,11),
TO_SIGNED(535,11),
TO_SIGNED(501,11),
TO_SIGNED(465,11),
TO_SIGNED(427,11),
TO_SIGNED(387,11),
TO_SIGNED(346,11),
TO_SIGNED(304,11),
TO_SIGNED(261,11),
TO_SIGNED(216,11),
TO_SIGNED(171,11),
TO_SIGNED(124,11),
TO_SIGNED(78,11),
TO_SIGNED(31,11),
TO_SIGNED(-16,11),
TO_SIGNED(-63,11),
TO_SIGNED(-110,11),
TO_SIGNED(-156,11),
TO_SIGNED(-202,11),
TO_SIGNED(-246,11),
TO_SIGNED(-290,11),
TO_SIGNED(-333,11),
TO_SIGNED(-375,11),
TO_SIGNED(-415,11),
TO_SIGNED(-453,11),
TO_SIGNED(-489,11),
TO_SIGNED(-524,11),
TO_SIGNED(-557,11),
TO_SIGNED(-587,11),
TO_SIGNED(-615,11),
TO_SIGNED(-641,11),
TO_SIGNED(-664,11),
TO_SIGNED(-685,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-730,11),
TO_SIGNED(-739,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-693,11),
TO_SIGNED(-673,11),
TO_SIGNED(-651,11),
TO_SIGNED(-627,11),
TO_SIGNED(-599,11),
TO_SIGNED(-570,11),
TO_SIGNED(-538,11),
TO_SIGNED(-505,11),
TO_SIGNED(-469,11),
TO_SIGNED(-431,11),
TO_SIGNED(-392,11),
TO_SIGNED(-351,11),
TO_SIGNED(-309,11),
TO_SIGNED(-266,11),
TO_SIGNED(-221,11),
TO_SIGNED(-176,11),
TO_SIGNED(-130,11),
TO_SIGNED(-83,11),
TO_SIGNED(-36,11),
TO_SIGNED(11,11),
TO_SIGNED(58,11),
TO_SIGNED(104,11),
TO_SIGNED(151,11),
TO_SIGNED(196,11),
TO_SIGNED(241,11),
TO_SIGNED(285,11),
TO_SIGNED(328,11),
TO_SIGNED(370,11),
TO_SIGNED(410,11),
TO_SIGNED(449,11),
TO_SIGNED(485,11),
TO_SIGNED(520,11),
TO_SIGNED(553,11),
TO_SIGNED(584,11),
TO_SIGNED(612,11),
TO_SIGNED(638,11),
TO_SIGNED(661,11),
TO_SIGNED(682,11),
TO_SIGNED(700,11),
TO_SIGNED(716,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(725,11),
TO_SIGNED(711,11),
TO_SIGNED(695,11),
TO_SIGNED(675,11),
TO_SIGNED(654,11),
TO_SIGNED(629,11),
TO_SIGNED(603,11),
TO_SIGNED(574,11),
TO_SIGNED(542,11),
TO_SIGNED(509,11),
TO_SIGNED(473,11),
TO_SIGNED(436,11),
TO_SIGNED(397,11),
TO_SIGNED(356,11),
TO_SIGNED(314,11),
TO_SIGNED(271,11),
TO_SIGNED(226,11),
TO_SIGNED(181,11),
TO_SIGNED(135,11),
TO_SIGNED(88,11),
TO_SIGNED(42,11),
TO_SIGNED(-5,11),
TO_SIGNED(-52,11),
TO_SIGNED(-99,11),
TO_SIGNED(-145,11),
TO_SIGNED(-191,11),
TO_SIGNED(-236,11),
TO_SIGNED(-280,11),
TO_SIGNED(-323,11),
TO_SIGNED(-365,11),
TO_SIGNED(-406,11),
TO_SIGNED(-444,11),
TO_SIGNED(-481,11),
TO_SIGNED(-516,11),
TO_SIGNED(-549,11),
TO_SIGNED(-580,11),
TO_SIGNED(-609,11),
TO_SIGNED(-635,11),
TO_SIGNED(-659,11),
TO_SIGNED(-680,11),
TO_SIGNED(-699,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-736,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-678,11),
TO_SIGNED(-656,11),
TO_SIGNED(-632,11),
TO_SIGNED(-606,11),
TO_SIGNED(-577,11),
TO_SIGNED(-546,11),
TO_SIGNED(-512,11),
TO_SIGNED(-477,11),
TO_SIGNED(-440,11),
TO_SIGNED(-401,11),
TO_SIGNED(-361,11),
TO_SIGNED(-319,11),
TO_SIGNED(-275,11),
TO_SIGNED(-231,11),
TO_SIGNED(-186,11),
TO_SIGNED(-140,11),
TO_SIGNED(-94,11),
TO_SIGNED(-47,11),
TO_SIGNED(0,11),
TO_SIGNED(47,11),
TO_SIGNED(94,11),
TO_SIGNED(140,11),
TO_SIGNED(186,11),
TO_SIGNED(231,11),
TO_SIGNED(275,11),
TO_SIGNED(319,11),
TO_SIGNED(361,11),
TO_SIGNED(401,11),
TO_SIGNED(440,11),
TO_SIGNED(477,11),
TO_SIGNED(512,11),
TO_SIGNED(546,11),
TO_SIGNED(577,11),
TO_SIGNED(606,11),
TO_SIGNED(632,11),
TO_SIGNED(656,11),
TO_SIGNED(678,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(736,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(699,11),
TO_SIGNED(680,11),
TO_SIGNED(659,11),
TO_SIGNED(635,11),
TO_SIGNED(609,11),
TO_SIGNED(580,11),
TO_SIGNED(549,11),
TO_SIGNED(516,11),
TO_SIGNED(481,11),
TO_SIGNED(444,11),
TO_SIGNED(406,11),
TO_SIGNED(365,11),
TO_SIGNED(323,11),
TO_SIGNED(280,11),
TO_SIGNED(236,11),
TO_SIGNED(191,11),
TO_SIGNED(145,11),
TO_SIGNED(99,11),
TO_SIGNED(52,11),
TO_SIGNED(5,11),
TO_SIGNED(-42,11),
TO_SIGNED(-88,11),
TO_SIGNED(-135,11),
TO_SIGNED(-181,11),
TO_SIGNED(-226,11),
TO_SIGNED(-271,11),
TO_SIGNED(-314,11),
TO_SIGNED(-356,11),
TO_SIGNED(-397,11),
TO_SIGNED(-436,11),
TO_SIGNED(-473,11),
TO_SIGNED(-509,11),
TO_SIGNED(-542,11),
TO_SIGNED(-574,11),
TO_SIGNED(-603,11),
TO_SIGNED(-629,11),
TO_SIGNED(-654,11),
TO_SIGNED(-675,11),
TO_SIGNED(-695,11),
TO_SIGNED(-711,11),
TO_SIGNED(-725,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-716,11),
TO_SIGNED(-700,11),
TO_SIGNED(-682,11),
TO_SIGNED(-661,11),
TO_SIGNED(-638,11),
TO_SIGNED(-612,11),
TO_SIGNED(-584,11),
TO_SIGNED(-553,11),
TO_SIGNED(-520,11),
TO_SIGNED(-485,11),
TO_SIGNED(-449,11),
TO_SIGNED(-410,11),
TO_SIGNED(-370,11),
TO_SIGNED(-328,11),
TO_SIGNED(-285,11),
TO_SIGNED(-241,11),
TO_SIGNED(-196,11),
TO_SIGNED(-151,11),
TO_SIGNED(-104,11),
TO_SIGNED(-58,11),
TO_SIGNED(-11,11),
TO_SIGNED(36,11),
TO_SIGNED(83,11),
TO_SIGNED(130,11),
TO_SIGNED(176,11),
TO_SIGNED(221,11),
TO_SIGNED(266,11),
TO_SIGNED(309,11),
TO_SIGNED(351,11),
TO_SIGNED(392,11),
TO_SIGNED(431,11),
TO_SIGNED(469,11),
TO_SIGNED(505,11),
TO_SIGNED(538,11),
TO_SIGNED(570,11),
TO_SIGNED(599,11),
TO_SIGNED(627,11),
TO_SIGNED(651,11),
TO_SIGNED(673,11),
TO_SIGNED(693,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(739,11),
TO_SIGNED(730,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(685,11),
TO_SIGNED(664,11),
TO_SIGNED(641,11),
TO_SIGNED(615,11),
TO_SIGNED(587,11),
TO_SIGNED(557,11),
TO_SIGNED(524,11),
TO_SIGNED(489,11),
TO_SIGNED(453,11),
TO_SIGNED(415,11),
TO_SIGNED(375,11),
TO_SIGNED(333,11),
TO_SIGNED(290,11),
TO_SIGNED(246,11),
TO_SIGNED(202,11),
TO_SIGNED(156,11),
TO_SIGNED(110,11),
TO_SIGNED(63,11),
TO_SIGNED(16,11),
TO_SIGNED(-31,11),
TO_SIGNED(-78,11),
TO_SIGNED(-124,11),
TO_SIGNED(-171,11),
TO_SIGNED(-216,11),
TO_SIGNED(-261,11),
TO_SIGNED(-304,11),
TO_SIGNED(-346,11),
TO_SIGNED(-387,11),
TO_SIGNED(-427,11),
TO_SIGNED(-465,11),
TO_SIGNED(-501,11),
TO_SIGNED(-535,11),
TO_SIGNED(-567,11),
TO_SIGNED(-596,11),
TO_SIGNED(-624,11),
TO_SIGNED(-648,11),
TO_SIGNED(-671,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-719,11),
TO_SIGNED(-704,11),
TO_SIGNED(-687,11),
TO_SIGNED(-666,11),
TO_SIGNED(-644,11),
TO_SIGNED(-618,11),
TO_SIGNED(-590,11),
TO_SIGNED(-560,11),
TO_SIGNED(-528,11),
TO_SIGNED(-493,11),
TO_SIGNED(-457,11),
TO_SIGNED(-419,11),
TO_SIGNED(-379,11),
TO_SIGNED(-338,11),
TO_SIGNED(-295,11),
TO_SIGNED(-251,11),
TO_SIGNED(-207,11),
TO_SIGNED(-161,11),
TO_SIGNED(-115,11),
TO_SIGNED(-68,11),
TO_SIGNED(-21,11),
TO_SIGNED(26,11),
TO_SIGNED(73,11),
TO_SIGNED(119,11),
TO_SIGNED(165,11),
TO_SIGNED(211,11),
TO_SIGNED(256,11),
TO_SIGNED(299,11),
TO_SIGNED(342,11),
TO_SIGNED(383,11),
TO_SIGNED(422,11),
TO_SIGNED(460,11),
TO_SIGNED(497,11),
TO_SIGNED(531,11),
TO_SIGNED(563,11),
TO_SIGNED(593,11),
TO_SIGNED(621,11),
TO_SIGNED(646,11),
TO_SIGNED(668,11),
TO_SIGNED(688,11),
TO_SIGNED(706,11),
TO_SIGNED(720,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(721,11),
TO_SIGNED(706,11),
TO_SIGNED(689,11),
TO_SIGNED(669,11),
TO_SIGNED(646,11),
TO_SIGNED(621,11),
TO_SIGNED(594,11),
TO_SIGNED(564,11),
TO_SIGNED(532,11),
TO_SIGNED(497,11),
TO_SIGNED(461,11),
TO_SIGNED(423,11),
TO_SIGNED(384,11),
TO_SIGNED(343,11),
TO_SIGNED(300,11),
TO_SIGNED(257,11),
TO_SIGNED(212,11),
TO_SIGNED(166,11),
TO_SIGNED(120,11),
TO_SIGNED(74,11),
TO_SIGNED(27,11),
TO_SIGNED(-20,11),
TO_SIGNED(-67,11),
TO_SIGNED(-114,11),
TO_SIGNED(-160,11),
TO_SIGNED(-206,11),
TO_SIGNED(-250,11),
TO_SIGNED(-294,11),
TO_SIGNED(-337,11),
TO_SIGNED(-378,11),
TO_SIGNED(-418,11),
TO_SIGNED(-456,11),
TO_SIGNED(-493,11),
TO_SIGNED(-527,11),
TO_SIGNED(-559,11),
TO_SIGNED(-590,11),
TO_SIGNED(-618,11),
TO_SIGNED(-643,11),
TO_SIGNED(-666,11),
TO_SIGNED(-686,11),
TO_SIGNED(-704,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-733,11),
TO_SIGNED(-722,11),
TO_SIGNED(-708,11),
TO_SIGNED(-691,11),
TO_SIGNED(-671,11),
TO_SIGNED(-649,11),
TO_SIGNED(-624,11),
TO_SIGNED(-597,11),
TO_SIGNED(-567,11),
TO_SIGNED(-535,11),
TO_SIGNED(-501,11),
TO_SIGNED(-466,11),
TO_SIGNED(-428,11),
TO_SIGNED(-388,11),
TO_SIGNED(-347,11),
TO_SIGNED(-305,11),
TO_SIGNED(-262,11),
TO_SIGNED(-217,11),
TO_SIGNED(-172,11),
TO_SIGNED(-125,11),
TO_SIGNED(-79,11),
TO_SIGNED(-32,11),
TO_SIGNED(15,11),
TO_SIGNED(62,11),
TO_SIGNED(109,11),
TO_SIGNED(155,11),
TO_SIGNED(201,11),
TO_SIGNED(245,11),
TO_SIGNED(289,11),
TO_SIGNED(332,11),
TO_SIGNED(374,11),
TO_SIGNED(414,11),
TO_SIGNED(452,11),
TO_SIGNED(489,11),
TO_SIGNED(523,11),
TO_SIGNED(556,11),
TO_SIGNED(586,11),
TO_SIGNED(615,11),
TO_SIGNED(640,11),
TO_SIGNED(663,11),
TO_SIGNED(684,11),
TO_SIGNED(702,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(710,11),
TO_SIGNED(693,11),
TO_SIGNED(674,11),
TO_SIGNED(652,11),
TO_SIGNED(627,11),
TO_SIGNED(600,11),
TO_SIGNED(571,11),
TO_SIGNED(539,11),
TO_SIGNED(505,11),
TO_SIGNED(470,11),
TO_SIGNED(432,11),
TO_SIGNED(393,11),
TO_SIGNED(352,11),
TO_SIGNED(310,11),
TO_SIGNED(267,11),
TO_SIGNED(222,11),
TO_SIGNED(177,11),
TO_SIGNED(131,11),
TO_SIGNED(84,11),
TO_SIGNED(37,11),
TO_SIGNED(-10,11),
TO_SIGNED(-57,11),
TO_SIGNED(-103,11),
TO_SIGNED(-150,11),
TO_SIGNED(-195,11),
TO_SIGNED(-240,11),
TO_SIGNED(-284,11),
TO_SIGNED(-327,11),
TO_SIGNED(-369,11),
TO_SIGNED(-409,11),
TO_SIGNED(-448,11),
TO_SIGNED(-485,11),
TO_SIGNED(-519,11),
TO_SIGNED(-552,11),
TO_SIGNED(-583,11),
TO_SIGNED(-611,11),
TO_SIGNED(-637,11),
TO_SIGNED(-661,11),
TO_SIGNED(-682,11),
TO_SIGNED(-700,11),
TO_SIGNED(-716,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-725,11),
TO_SIGNED(-711,11),
TO_SIGNED(-695,11),
TO_SIGNED(-676,11),
TO_SIGNED(-654,11),
TO_SIGNED(-630,11),
TO_SIGNED(-603,11),
TO_SIGNED(-574,11),
TO_SIGNED(-543,11),
TO_SIGNED(-509,11),
TO_SIGNED(-474,11),
TO_SIGNED(-437,11),
TO_SIGNED(-397,11),
TO_SIGNED(-357,11),
TO_SIGNED(-315,11),
TO_SIGNED(-272,11),
TO_SIGNED(-227,11),
TO_SIGNED(-182,11),
TO_SIGNED(-136,11),
TO_SIGNED(-90,11),
TO_SIGNED(-43,11),
TO_SIGNED(4,11),
TO_SIGNED(51,11),
TO_SIGNED(98,11),
TO_SIGNED(144,11),
TO_SIGNED(190,11),
TO_SIGNED(235,11),
TO_SIGNED(279,11),
TO_SIGNED(323,11),
TO_SIGNED(364,11),
TO_SIGNED(405,11),
TO_SIGNED(443,11),
TO_SIGNED(480,11),
TO_SIGNED(516,11),
TO_SIGNED(549,11),
TO_SIGNED(580,11),
TO_SIGNED(608,11),
TO_SIGNED(635,11),
TO_SIGNED(658,11),
TO_SIGNED(680,11),
TO_SIGNED(698,11),
TO_SIGNED(714,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(713,11),
TO_SIGNED(697,11),
TO_SIGNED(678,11),
TO_SIGNED(657,11),
TO_SIGNED(633,11),
TO_SIGNED(606,11),
TO_SIGNED(578,11),
TO_SIGNED(547,11),
TO_SIGNED(513,11),
TO_SIGNED(478,11),
TO_SIGNED(441,11),
TO_SIGNED(402,11),
TO_SIGNED(362,11),
TO_SIGNED(320,11),
TO_SIGNED(276,11),
TO_SIGNED(232,11),
TO_SIGNED(187,11),
TO_SIGNED(141,11),
TO_SIGNED(95,11),
TO_SIGNED(48,11),
TO_SIGNED(1,11),
TO_SIGNED(-46,11),
TO_SIGNED(-93,11),
TO_SIGNED(-139,11),
TO_SIGNED(-185,11),
TO_SIGNED(-230,11),
TO_SIGNED(-275,11),
TO_SIGNED(-318,11),
TO_SIGNED(-360,11),
TO_SIGNED(-400,11),
TO_SIGNED(-439,11),
TO_SIGNED(-476,11),
TO_SIGNED(-512,11),
TO_SIGNED(-545,11),
TO_SIGNED(-576,11),
TO_SIGNED(-605,11),
TO_SIGNED(-632,11),
TO_SIGNED(-656,11),
TO_SIGNED(-677,11),
TO_SIGNED(-696,11),
TO_SIGNED(-712,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-715,11),
TO_SIGNED(-699,11),
TO_SIGNED(-681,11),
TO_SIGNED(-659,11),
TO_SIGNED(-636,11),
TO_SIGNED(-610,11),
TO_SIGNED(-581,11),
TO_SIGNED(-550,11),
TO_SIGNED(-517,11),
TO_SIGNED(-482,11),
TO_SIGNED(-445,11),
TO_SIGNED(-406,11),
TO_SIGNED(-366,11),
TO_SIGNED(-324,11),
TO_SIGNED(-281,11),
TO_SIGNED(-237,11),
TO_SIGNED(-192,11),
TO_SIGNED(-147,11),
TO_SIGNED(-100,11),
TO_SIGNED(-53,11),
TO_SIGNED(-6,11),
TO_SIGNED(41,11),
TO_SIGNED(87,11),
TO_SIGNED(134,11),
TO_SIGNED(180,11),
TO_SIGNED(225,11),
TO_SIGNED(270,11),
TO_SIGNED(313,11),
TO_SIGNED(355,11),
TO_SIGNED(396,11),
TO_SIGNED(435,11),
TO_SIGNED(472,11),
TO_SIGNED(508,11),
TO_SIGNED(541,11),
TO_SIGNED(573,11),
TO_SIGNED(602,11),
TO_SIGNED(629,11),
TO_SIGNED(653,11),
TO_SIGNED(675,11),
TO_SIGNED(694,11),
TO_SIGNED(711,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(729,11),
TO_SIGNED(716,11),
TO_SIGNED(701,11),
TO_SIGNED(683,11),
TO_SIGNED(662,11),
TO_SIGNED(639,11),
TO_SIGNED(613,11),
TO_SIGNED(584,11),
TO_SIGNED(554,11),
TO_SIGNED(521,11),
TO_SIGNED(486,11),
TO_SIGNED(449,11),
TO_SIGNED(411,11),
TO_SIGNED(371,11),
TO_SIGNED(329,11),
TO_SIGNED(286,11),
TO_SIGNED(242,11),
TO_SIGNED(197,11),
TO_SIGNED(152,11),
TO_SIGNED(105,11),
TO_SIGNED(59,11),
TO_SIGNED(12,11),
TO_SIGNED(-35,11),
TO_SIGNED(-82,11),
TO_SIGNED(-129,11),
TO_SIGNED(-175,11),
TO_SIGNED(-220,11),
TO_SIGNED(-265,11),
TO_SIGNED(-308,11),
TO_SIGNED(-350,11),
TO_SIGNED(-391,11),
TO_SIGNED(-430,11),
TO_SIGNED(-468,11),
TO_SIGNED(-504,11),
TO_SIGNED(-538,11),
TO_SIGNED(-569,11),
TO_SIGNED(-599,11),
TO_SIGNED(-626,11),
TO_SIGNED(-651,11),
TO_SIGNED(-673,11),
TO_SIGNED(-692,11),
TO_SIGNED(-709,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-685,11),
TO_SIGNED(-664,11),
TO_SIGNED(-641,11),
TO_SIGNED(-616,11),
TO_SIGNED(-588,11),
TO_SIGNED(-557,11),
TO_SIGNED(-525,11),
TO_SIGNED(-490,11),
TO_SIGNED(-454,11),
TO_SIGNED(-415,11),
TO_SIGNED(-375,11),
TO_SIGNED(-334,11),
TO_SIGNED(-291,11),
TO_SIGNED(-247,11),
TO_SIGNED(-203,11),
TO_SIGNED(-157,11),
TO_SIGNED(-111,11),
TO_SIGNED(-64,11),
TO_SIGNED(-17,11),
TO_SIGNED(30,11),
TO_SIGNED(77,11),
TO_SIGNED(123,11),
TO_SIGNED(169,11),
TO_SIGNED(215,11),
TO_SIGNED(260,11),
TO_SIGNED(303,11),
TO_SIGNED(345,11),
TO_SIGNED(387,11),
TO_SIGNED(426,11),
TO_SIGNED(464,11),
TO_SIGNED(500,11),
TO_SIGNED(534,11),
TO_SIGNED(566,11),
TO_SIGNED(596,11),
TO_SIGNED(623,11),
TO_SIGNED(648,11),
TO_SIGNED(670,11),
TO_SIGNED(690,11),
TO_SIGNED(707,11),
TO_SIGNED(721,11),
TO_SIGNED(733,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(705,11),
TO_SIGNED(687,11),
TO_SIGNED(667,11),
TO_SIGNED(644,11),
TO_SIGNED(619,11),
TO_SIGNED(591,11),
TO_SIGNED(561,11),
TO_SIGNED(529,11),
TO_SIGNED(494,11),
TO_SIGNED(458,11),
TO_SIGNED(420,11),
TO_SIGNED(380,11),
TO_SIGNED(339,11),
TO_SIGNED(296,11),
TO_SIGNED(252,11),
TO_SIGNED(208,11),
TO_SIGNED(162,11),
TO_SIGNED(116,11),
TO_SIGNED(69,11),
TO_SIGNED(22,11),
TO_SIGNED(-25,11),
TO_SIGNED(-71,11),
TO_SIGNED(-118,11),
TO_SIGNED(-164,11),
TO_SIGNED(-210,11),
TO_SIGNED(-255,11),
TO_SIGNED(-298,11),
TO_SIGNED(-341,11),
TO_SIGNED(-382,11),
TO_SIGNED(-422,11),
TO_SIGNED(-460,11),
TO_SIGNED(-496,11),
TO_SIGNED(-530,11),
TO_SIGNED(-562,11),
TO_SIGNED(-592,11),
TO_SIGNED(-620,11),
TO_SIGNED(-645,11),
TO_SIGNED(-668,11),
TO_SIGNED(-688,11),
TO_SIGNED(-705,11),
TO_SIGNED(-720,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-721,11),
TO_SIGNED(-706,11),
TO_SIGNED(-689,11),
TO_SIGNED(-669,11),
TO_SIGNED(-647,11),
TO_SIGNED(-622,11),
TO_SIGNED(-594,11),
TO_SIGNED(-564,11),
TO_SIGNED(-532,11),
TO_SIGNED(-498,11),
TO_SIGNED(-462,11),
TO_SIGNED(-424,11),
TO_SIGNED(-385,11),
TO_SIGNED(-344,11),
TO_SIGNED(-301,11),
TO_SIGNED(-258,11),
TO_SIGNED(-213,11),
TO_SIGNED(-167,11),
TO_SIGNED(-121,11),
TO_SIGNED(-75,11),
TO_SIGNED(-28,11),
TO_SIGNED(19,11),
TO_SIGNED(66,11),
TO_SIGNED(113,11),
TO_SIGNED(159,11),
TO_SIGNED(205,11),
TO_SIGNED(249,11),
TO_SIGNED(293,11),
TO_SIGNED(336,11),
TO_SIGNED(377,11),
TO_SIGNED(417,11),
TO_SIGNED(455,11),
TO_SIGNED(492,11),
TO_SIGNED(526,11),
TO_SIGNED(559,11),
TO_SIGNED(589,11),
TO_SIGNED(617,11),
TO_SIGNED(642,11),
TO_SIGNED(665,11),
TO_SIGNED(686,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(708,11),
TO_SIGNED(691,11),
TO_SIGNED(672,11),
TO_SIGNED(650,11),
TO_SIGNED(625,11),
TO_SIGNED(598,11),
TO_SIGNED(568,11),
TO_SIGNED(536,11),
TO_SIGNED(502,11),
TO_SIGNED(466,11),
TO_SIGNED(429,11),
TO_SIGNED(389,11),
TO_SIGNED(348,11),
TO_SIGNED(306,11),
TO_SIGNED(263,11),
TO_SIGNED(218,11),
TO_SIGNED(173,11),
TO_SIGNED(127,11),
TO_SIGNED(80,11),
TO_SIGNED(33,11),
TO_SIGNED(-14,11),
TO_SIGNED(-61,11),
TO_SIGNED(-108,11),
TO_SIGNED(-154,11),
TO_SIGNED(-200,11),
TO_SIGNED(-244,11),
TO_SIGNED(-288,11),
TO_SIGNED(-331,11),
TO_SIGNED(-373,11),
TO_SIGNED(-413,11),
TO_SIGNED(-451,11),
TO_SIGNED(-488,11),
TO_SIGNED(-523,11),
TO_SIGNED(-555,11),
TO_SIGNED(-586,11),
TO_SIGNED(-614,11),
TO_SIGNED(-640,11),
TO_SIGNED(-663,11),
TO_SIGNED(-684,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-729,11),
TO_SIGNED(-739,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-710,11),
TO_SIGNED(-693,11),
TO_SIGNED(-674,11),
TO_SIGNED(-652,11),
TO_SIGNED(-628,11),
TO_SIGNED(-601,11),
TO_SIGNED(-571,11),
TO_SIGNED(-540,11),
TO_SIGNED(-506,11),
TO_SIGNED(-471,11),
TO_SIGNED(-433,11),
TO_SIGNED(-394,11),
TO_SIGNED(-353,11),
TO_SIGNED(-311,11),
TO_SIGNED(-268,11),
TO_SIGNED(-223,11),
TO_SIGNED(-178,11),
TO_SIGNED(-132,11),
TO_SIGNED(-85,11),
TO_SIGNED(-38,11),
TO_SIGNED(9,11),
TO_SIGNED(56,11),
TO_SIGNED(102,11),
TO_SIGNED(149,11),
TO_SIGNED(194,11),
TO_SIGNED(239,11),
TO_SIGNED(283,11),
TO_SIGNED(326,11),
TO_SIGNED(368,11),
TO_SIGNED(408,11),
TO_SIGNED(447,11),
TO_SIGNED(484,11),
TO_SIGNED(519,11),
TO_SIGNED(552,11),
TO_SIGNED(582,11),
TO_SIGNED(611,11),
TO_SIGNED(637,11),
TO_SIGNED(660,11),
TO_SIGNED(681,11),
TO_SIGNED(700,11),
TO_SIGNED(715,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(736,11),
TO_SIGNED(725,11),
TO_SIGNED(712,11),
TO_SIGNED(695,11),
TO_SIGNED(676,11),
TO_SIGNED(655,11),
TO_SIGNED(631,11),
TO_SIGNED(604,11),
TO_SIGNED(575,11),
TO_SIGNED(544,11),
TO_SIGNED(510,11),
TO_SIGNED(475,11),
TO_SIGNED(437,11),
TO_SIGNED(398,11),
TO_SIGNED(358,11),
TO_SIGNED(316,11),
TO_SIGNED(273,11),
TO_SIGNED(228,11),
TO_SIGNED(183,11),
TO_SIGNED(137,11),
TO_SIGNED(91,11),
TO_SIGNED(44,11),
TO_SIGNED(-3,11),
TO_SIGNED(-50,11),
TO_SIGNED(-97,11),
TO_SIGNED(-143,11),
TO_SIGNED(-189,11),
TO_SIGNED(-234,11),
TO_SIGNED(-278,11),
TO_SIGNED(-322,11),
TO_SIGNED(-363,11),
TO_SIGNED(-404,11),
TO_SIGNED(-443,11),
TO_SIGNED(-480,11),
TO_SIGNED(-515,11),
TO_SIGNED(-548,11),
TO_SIGNED(-579,11),
TO_SIGNED(-608,11),
TO_SIGNED(-634,11),
TO_SIGNED(-658,11),
TO_SIGNED(-679,11),
TO_SIGNED(-698,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-679,11),
TO_SIGNED(-657,11),
TO_SIGNED(-633,11),
TO_SIGNED(-607,11),
TO_SIGNED(-578,11),
TO_SIGNED(-547,11),
TO_SIGNED(-514,11),
TO_SIGNED(-479,11),
TO_SIGNED(-442,11),
TO_SIGNED(-403,11),
TO_SIGNED(-362,11),
TO_SIGNED(-321,11),
TO_SIGNED(-277,11),
TO_SIGNED(-233,11),
TO_SIGNED(-188,11),
TO_SIGNED(-142,11),
TO_SIGNED(-96,11),
TO_SIGNED(-49,11),
TO_SIGNED(-2,11),
TO_SIGNED(45,11),
TO_SIGNED(92,11),
TO_SIGNED(138,11),
TO_SIGNED(184,11),
TO_SIGNED(229,11),
TO_SIGNED(274,11),
TO_SIGNED(317,11),
TO_SIGNED(359,11),
TO_SIGNED(399,11),
TO_SIGNED(438,11),
TO_SIGNED(476,11),
TO_SIGNED(511,11),
TO_SIGNED(544,11),
TO_SIGNED(576,11),
TO_SIGNED(605,11),
TO_SIGNED(631,11),
TO_SIGNED(655,11),
TO_SIGNED(677,11),
TO_SIGNED(696,11),
TO_SIGNED(712,11),
TO_SIGNED(725,11),
TO_SIGNED(736,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(715,11),
TO_SIGNED(699,11),
TO_SIGNED(681,11),
TO_SIGNED(660,11),
TO_SIGNED(636,11),
TO_SIGNED(610,11),
TO_SIGNED(582,11),
TO_SIGNED(551,11),
TO_SIGNED(518,11),
TO_SIGNED(483,11),
TO_SIGNED(446,11),
TO_SIGNED(407,11),
TO_SIGNED(367,11),
TO_SIGNED(325,11),
TO_SIGNED(282,11),
TO_SIGNED(238,11),
TO_SIGNED(193,11),
TO_SIGNED(148,11),
TO_SIGNED(101,11),
TO_SIGNED(54,11),
TO_SIGNED(7,11),
TO_SIGNED(-40,11),
TO_SIGNED(-86,11),
TO_SIGNED(-133,11),
TO_SIGNED(-179,11),
TO_SIGNED(-224,11),
TO_SIGNED(-269,11),
TO_SIGNED(-312,11),
TO_SIGNED(-354,11),
TO_SIGNED(-395,11),
TO_SIGNED(-434,11),
TO_SIGNED(-471,11),
TO_SIGNED(-507,11),
TO_SIGNED(-541,11),
TO_SIGNED(-572,11),
TO_SIGNED(-601,11),
TO_SIGNED(-628,11),
TO_SIGNED(-653,11),
TO_SIGNED(-675,11),
TO_SIGNED(-694,11),
TO_SIGNED(-710,11),
TO_SIGNED(-724,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-701,11),
TO_SIGNED(-683,11),
TO_SIGNED(-662,11),
TO_SIGNED(-639,11),
TO_SIGNED(-613,11),
TO_SIGNED(-585,11),
TO_SIGNED(-554,11),
TO_SIGNED(-522,11),
TO_SIGNED(-487,11),
TO_SIGNED(-450,11),
TO_SIGNED(-412,11),
TO_SIGNED(-372,11),
TO_SIGNED(-330,11),
TO_SIGNED(-287,11),
TO_SIGNED(-243,11),
TO_SIGNED(-198,11),
TO_SIGNED(-153,11),
TO_SIGNED(-106,11),
TO_SIGNED(-60,11),
TO_SIGNED(-13,11),
TO_SIGNED(34,11),
TO_SIGNED(81,11),
TO_SIGNED(128,11),
TO_SIGNED(174,11),
TO_SIGNED(219,11),
TO_SIGNED(264,11),
TO_SIGNED(307,11),
TO_SIGNED(349,11),
TO_SIGNED(390,11),
TO_SIGNED(430,11),
TO_SIGNED(467,11),
TO_SIGNED(503,11),
TO_SIGNED(537,11),
TO_SIGNED(569,11),
TO_SIGNED(598,11),
TO_SIGNED(625,11),
TO_SIGNED(650,11),
TO_SIGNED(672,11),
TO_SIGNED(692,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(730,11),
TO_SIGNED(718,11),
TO_SIGNED(703,11),
TO_SIGNED(685,11),
TO_SIGNED(665,11),
TO_SIGNED(642,11),
TO_SIGNED(616,11),
TO_SIGNED(588,11),
TO_SIGNED(558,11),
TO_SIGNED(526,11),
TO_SIGNED(491,11),
TO_SIGNED(455,11),
TO_SIGNED(416,11),
TO_SIGNED(376,11),
TO_SIGNED(335,11),
TO_SIGNED(292,11),
TO_SIGNED(248,11),
TO_SIGNED(204,11),
TO_SIGNED(158,11),
TO_SIGNED(112,11),
TO_SIGNED(65,11),
TO_SIGNED(18,11),
TO_SIGNED(-29,11),
TO_SIGNED(-76,11),
TO_SIGNED(-122,11),
TO_SIGNED(-168,11),
TO_SIGNED(-214,11),
TO_SIGNED(-259,11),
TO_SIGNED(-302,11),
TO_SIGNED(-345,11),
TO_SIGNED(-386,11),
TO_SIGNED(-425,11),
TO_SIGNED(-463,11),
TO_SIGNED(-499,11),
TO_SIGNED(-533,11),
TO_SIGNED(-565,11),
TO_SIGNED(-595,11),
TO_SIGNED(-622,11),
TO_SIGNED(-647,11),
TO_SIGNED(-670,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-721,11),
TO_SIGNED(-733,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-720,11),
TO_SIGNED(-705,11),
TO_SIGNED(-688,11),
TO_SIGNED(-667,11),
TO_SIGNED(-645,11),
TO_SIGNED(-619,11),
TO_SIGNED(-592,11),
TO_SIGNED(-562,11),
TO_SIGNED(-529,11),
TO_SIGNED(-495,11),
TO_SIGNED(-459,11),
TO_SIGNED(-421,11),
TO_SIGNED(-381,11),
TO_SIGNED(-340,11),
TO_SIGNED(-297,11),
TO_SIGNED(-254,11),
TO_SIGNED(-209,11),
TO_SIGNED(-163,11),
TO_SIGNED(-117,11),
TO_SIGNED(-70,11),
TO_SIGNED(-24,11),
TO_SIGNED(24,11),
TO_SIGNED(70,11),
TO_SIGNED(117,11),
TO_SIGNED(163,11),
TO_SIGNED(209,11),
TO_SIGNED(254,11),
TO_SIGNED(297,11),
TO_SIGNED(340,11),
TO_SIGNED(381,11),
TO_SIGNED(421,11),
TO_SIGNED(459,11),
TO_SIGNED(495,11),
TO_SIGNED(529,11),
TO_SIGNED(562,11),
TO_SIGNED(592,11),
TO_SIGNED(619,11),
TO_SIGNED(645,11),
TO_SIGNED(667,11),
TO_SIGNED(688,11),
TO_SIGNED(705,11),
TO_SIGNED(720,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(733,11),
TO_SIGNED(721,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(670,11),
TO_SIGNED(647,11),
TO_SIGNED(622,11),
TO_SIGNED(595,11),
TO_SIGNED(565,11),
TO_SIGNED(533,11),
TO_SIGNED(499,11),
TO_SIGNED(463,11),
TO_SIGNED(425,11),
TO_SIGNED(386,11),
TO_SIGNED(345,11),
TO_SIGNED(302,11),
TO_SIGNED(259,11),
TO_SIGNED(214,11),
TO_SIGNED(168,11),
TO_SIGNED(122,11),
TO_SIGNED(76,11),
TO_SIGNED(29,11),
TO_SIGNED(-18,11),
TO_SIGNED(-65,11),
TO_SIGNED(-112,11),
TO_SIGNED(-158,11),
TO_SIGNED(-204,11),
TO_SIGNED(-248,11),
TO_SIGNED(-292,11),
TO_SIGNED(-335,11),
TO_SIGNED(-376,11),
TO_SIGNED(-416,11),
TO_SIGNED(-455,11),
TO_SIGNED(-491,11),
TO_SIGNED(-526,11),
TO_SIGNED(-558,11),
TO_SIGNED(-588,11),
TO_SIGNED(-616,11),
TO_SIGNED(-642,11),
TO_SIGNED(-665,11),
TO_SIGNED(-685,11),
TO_SIGNED(-703,11),
TO_SIGNED(-718,11),
TO_SIGNED(-730,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-692,11),
TO_SIGNED(-672,11),
TO_SIGNED(-650,11),
TO_SIGNED(-625,11),
TO_SIGNED(-598,11),
TO_SIGNED(-569,11),
TO_SIGNED(-537,11),
TO_SIGNED(-503,11),
TO_SIGNED(-467,11),
TO_SIGNED(-430,11),
TO_SIGNED(-390,11),
TO_SIGNED(-349,11),
TO_SIGNED(-307,11),
TO_SIGNED(-264,11),
TO_SIGNED(-219,11),
TO_SIGNED(-174,11),
TO_SIGNED(-128,11),
TO_SIGNED(-81,11),
TO_SIGNED(-34,11),
TO_SIGNED(13,11),
TO_SIGNED(60,11),
TO_SIGNED(106,11),
TO_SIGNED(153,11),
TO_SIGNED(198,11),
TO_SIGNED(243,11),
TO_SIGNED(287,11),
TO_SIGNED(330,11),
TO_SIGNED(372,11),
TO_SIGNED(412,11),
TO_SIGNED(450,11),
TO_SIGNED(487,11),
TO_SIGNED(522,11),
TO_SIGNED(554,11),
TO_SIGNED(585,11),
TO_SIGNED(613,11),
TO_SIGNED(639,11),
TO_SIGNED(662,11),
TO_SIGNED(683,11),
TO_SIGNED(701,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(724,11),
TO_SIGNED(710,11),
TO_SIGNED(694,11),
TO_SIGNED(675,11),
TO_SIGNED(653,11),
TO_SIGNED(628,11),
TO_SIGNED(601,11),
TO_SIGNED(572,11),
TO_SIGNED(541,11),
TO_SIGNED(507,11),
TO_SIGNED(471,11),
TO_SIGNED(434,11),
TO_SIGNED(395,11),
TO_SIGNED(354,11),
TO_SIGNED(312,11),
TO_SIGNED(269,11),
TO_SIGNED(224,11),
TO_SIGNED(179,11),
TO_SIGNED(133,11),
TO_SIGNED(86,11),
TO_SIGNED(40,11),
TO_SIGNED(-7,11),
TO_SIGNED(-54,11),
TO_SIGNED(-101,11),
TO_SIGNED(-148,11),
TO_SIGNED(-193,11),
TO_SIGNED(-238,11),
TO_SIGNED(-282,11),
TO_SIGNED(-325,11),
TO_SIGNED(-367,11),
TO_SIGNED(-407,11),
TO_SIGNED(-446,11),
TO_SIGNED(-483,11),
TO_SIGNED(-518,11),
TO_SIGNED(-551,11),
TO_SIGNED(-582,11),
TO_SIGNED(-610,11),
TO_SIGNED(-636,11),
TO_SIGNED(-660,11),
TO_SIGNED(-681,11),
TO_SIGNED(-699,11),
TO_SIGNED(-715,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-736,11),
TO_SIGNED(-725,11),
TO_SIGNED(-712,11),
TO_SIGNED(-696,11),
TO_SIGNED(-677,11),
TO_SIGNED(-655,11),
TO_SIGNED(-631,11),
TO_SIGNED(-605,11),
TO_SIGNED(-576,11),
TO_SIGNED(-544,11),
TO_SIGNED(-511,11),
TO_SIGNED(-476,11),
TO_SIGNED(-438,11),
TO_SIGNED(-399,11),
TO_SIGNED(-359,11),
TO_SIGNED(-317,11),
TO_SIGNED(-274,11),
TO_SIGNED(-229,11),
TO_SIGNED(-184,11),
TO_SIGNED(-138,11),
TO_SIGNED(-92,11),
TO_SIGNED(-45,11),
TO_SIGNED(2,11),
TO_SIGNED(49,11),
TO_SIGNED(96,11),
TO_SIGNED(142,11),
TO_SIGNED(188,11),
TO_SIGNED(233,11),
TO_SIGNED(277,11),
TO_SIGNED(321,11),
TO_SIGNED(362,11),
TO_SIGNED(403,11),
TO_SIGNED(442,11),
TO_SIGNED(479,11),
TO_SIGNED(514,11),
TO_SIGNED(547,11),
TO_SIGNED(578,11),
TO_SIGNED(607,11),
TO_SIGNED(633,11),
TO_SIGNED(657,11),
TO_SIGNED(679,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(698,11),
TO_SIGNED(679,11),
TO_SIGNED(658,11),
TO_SIGNED(634,11),
TO_SIGNED(608,11),
TO_SIGNED(579,11),
TO_SIGNED(548,11),
TO_SIGNED(515,11),
TO_SIGNED(480,11),
TO_SIGNED(443,11),
TO_SIGNED(404,11),
TO_SIGNED(363,11),
TO_SIGNED(322,11),
TO_SIGNED(278,11),
TO_SIGNED(234,11),
TO_SIGNED(189,11),
TO_SIGNED(143,11),
TO_SIGNED(97,11),
TO_SIGNED(50,11),
TO_SIGNED(3,11),
TO_SIGNED(-44,11),
TO_SIGNED(-91,11),
TO_SIGNED(-137,11),
TO_SIGNED(-183,11),
TO_SIGNED(-228,11),
TO_SIGNED(-273,11),
TO_SIGNED(-316,11),
TO_SIGNED(-358,11),
TO_SIGNED(-398,11),
TO_SIGNED(-437,11),
TO_SIGNED(-475,11),
TO_SIGNED(-510,11),
TO_SIGNED(-544,11),
TO_SIGNED(-575,11),
TO_SIGNED(-604,11),
TO_SIGNED(-631,11),
TO_SIGNED(-655,11),
TO_SIGNED(-676,11),
TO_SIGNED(-695,11),
TO_SIGNED(-712,11),
TO_SIGNED(-725,11),
TO_SIGNED(-736,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-715,11),
TO_SIGNED(-700,11),
TO_SIGNED(-681,11),
TO_SIGNED(-660,11),
TO_SIGNED(-637,11),
TO_SIGNED(-611,11),
TO_SIGNED(-582,11),
TO_SIGNED(-552,11),
TO_SIGNED(-519,11),
TO_SIGNED(-484,11),
TO_SIGNED(-447,11),
TO_SIGNED(-408,11),
TO_SIGNED(-368,11),
TO_SIGNED(-326,11),
TO_SIGNED(-283,11),
TO_SIGNED(-239,11),
TO_SIGNED(-194,11),
TO_SIGNED(-149,11),
TO_SIGNED(-102,11),
TO_SIGNED(-56,11),
TO_SIGNED(-9,11),
TO_SIGNED(38,11),
TO_SIGNED(85,11),
TO_SIGNED(132,11),
TO_SIGNED(178,11),
TO_SIGNED(223,11),
TO_SIGNED(268,11),
TO_SIGNED(311,11),
TO_SIGNED(353,11),
TO_SIGNED(394,11),
TO_SIGNED(433,11),
TO_SIGNED(471,11),
TO_SIGNED(506,11),
TO_SIGNED(540,11),
TO_SIGNED(571,11),
TO_SIGNED(601,11),
TO_SIGNED(628,11),
TO_SIGNED(652,11),
TO_SIGNED(674,11),
TO_SIGNED(693,11),
TO_SIGNED(710,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(739,11),
TO_SIGNED(729,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(684,11),
TO_SIGNED(663,11),
TO_SIGNED(640,11),
TO_SIGNED(614,11),
TO_SIGNED(586,11),
TO_SIGNED(555,11),
TO_SIGNED(523,11),
TO_SIGNED(488,11),
TO_SIGNED(451,11),
TO_SIGNED(413,11),
TO_SIGNED(373,11),
TO_SIGNED(331,11),
TO_SIGNED(288,11),
TO_SIGNED(244,11),
TO_SIGNED(200,11),
TO_SIGNED(154,11),
TO_SIGNED(108,11),
TO_SIGNED(61,11),
TO_SIGNED(14,11),
TO_SIGNED(-33,11),
TO_SIGNED(-80,11),
TO_SIGNED(-127,11),
TO_SIGNED(-173,11),
TO_SIGNED(-218,11),
TO_SIGNED(-263,11),
TO_SIGNED(-306,11),
TO_SIGNED(-348,11),
TO_SIGNED(-389,11),
TO_SIGNED(-429,11),
TO_SIGNED(-466,11),
TO_SIGNED(-502,11),
TO_SIGNED(-536,11),
TO_SIGNED(-568,11),
TO_SIGNED(-598,11),
TO_SIGNED(-625,11),
TO_SIGNED(-650,11),
TO_SIGNED(-672,11),
TO_SIGNED(-691,11),
TO_SIGNED(-708,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-686,11),
TO_SIGNED(-665,11),
TO_SIGNED(-642,11),
TO_SIGNED(-617,11),
TO_SIGNED(-589,11),
TO_SIGNED(-559,11),
TO_SIGNED(-526,11),
TO_SIGNED(-492,11),
TO_SIGNED(-455,11),
TO_SIGNED(-417,11),
TO_SIGNED(-377,11),
TO_SIGNED(-336,11),
TO_SIGNED(-293,11),
TO_SIGNED(-249,11),
TO_SIGNED(-205,11),
TO_SIGNED(-159,11),
TO_SIGNED(-113,11),
TO_SIGNED(-66,11),
TO_SIGNED(-19,11),
TO_SIGNED(28,11),
TO_SIGNED(75,11),
TO_SIGNED(121,11),
TO_SIGNED(167,11),
TO_SIGNED(213,11),
TO_SIGNED(258,11),
TO_SIGNED(301,11),
TO_SIGNED(344,11),
TO_SIGNED(385,11),
TO_SIGNED(424,11),
TO_SIGNED(462,11),
TO_SIGNED(498,11),
TO_SIGNED(532,11),
TO_SIGNED(564,11),
TO_SIGNED(594,11),
TO_SIGNED(622,11),
TO_SIGNED(647,11),
TO_SIGNED(669,11),
TO_SIGNED(689,11),
TO_SIGNED(706,11),
TO_SIGNED(721,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(720,11),
TO_SIGNED(705,11),
TO_SIGNED(688,11),
TO_SIGNED(668,11),
TO_SIGNED(645,11),
TO_SIGNED(620,11),
TO_SIGNED(592,11),
TO_SIGNED(562,11),
TO_SIGNED(530,11),
TO_SIGNED(496,11),
TO_SIGNED(460,11),
TO_SIGNED(422,11),
TO_SIGNED(382,11),
TO_SIGNED(341,11),
TO_SIGNED(298,11),
TO_SIGNED(255,11),
TO_SIGNED(210,11),
TO_SIGNED(164,11),
TO_SIGNED(118,11),
TO_SIGNED(71,11),
TO_SIGNED(25,11),
TO_SIGNED(-22,11),
TO_SIGNED(-69,11),
TO_SIGNED(-116,11),
TO_SIGNED(-162,11),
TO_SIGNED(-208,11),
TO_SIGNED(-252,11),
TO_SIGNED(-296,11),
TO_SIGNED(-339,11),
TO_SIGNED(-380,11),
TO_SIGNED(-420,11),
TO_SIGNED(-458,11),
TO_SIGNED(-494,11),
TO_SIGNED(-529,11),
TO_SIGNED(-561,11),
TO_SIGNED(-591,11),
TO_SIGNED(-619,11),
TO_SIGNED(-644,11),
TO_SIGNED(-667,11),
TO_SIGNED(-687,11),
TO_SIGNED(-705,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-733,11),
TO_SIGNED(-721,11),
TO_SIGNED(-707,11),
TO_SIGNED(-690,11),
TO_SIGNED(-670,11),
TO_SIGNED(-648,11),
TO_SIGNED(-623,11),
TO_SIGNED(-596,11),
TO_SIGNED(-566,11),
TO_SIGNED(-534,11),
TO_SIGNED(-500,11),
TO_SIGNED(-464,11),
TO_SIGNED(-426,11),
TO_SIGNED(-387,11),
TO_SIGNED(-345,11),
TO_SIGNED(-303,11),
TO_SIGNED(-260,11),
TO_SIGNED(-215,11),
TO_SIGNED(-169,11),
TO_SIGNED(-123,11),
TO_SIGNED(-77,11),
TO_SIGNED(-30,11),
TO_SIGNED(17,11),
TO_SIGNED(64,11),
TO_SIGNED(111,11),
TO_SIGNED(157,11),
TO_SIGNED(203,11),
TO_SIGNED(247,11),
TO_SIGNED(291,11),
TO_SIGNED(334,11),
TO_SIGNED(375,11),
TO_SIGNED(415,11),
TO_SIGNED(454,11),
TO_SIGNED(490,11),
TO_SIGNED(525,11),
TO_SIGNED(557,11),
TO_SIGNED(588,11),
TO_SIGNED(616,11),
TO_SIGNED(641,11),
TO_SIGNED(664,11),
TO_SIGNED(685,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(709,11),
TO_SIGNED(692,11),
TO_SIGNED(673,11),
TO_SIGNED(651,11),
TO_SIGNED(626,11),
TO_SIGNED(599,11),
TO_SIGNED(569,11),
TO_SIGNED(538,11),
TO_SIGNED(504,11),
TO_SIGNED(468,11),
TO_SIGNED(430,11),
TO_SIGNED(391,11),
TO_SIGNED(350,11),
TO_SIGNED(308,11),
TO_SIGNED(265,11),
TO_SIGNED(220,11),
TO_SIGNED(175,11),
TO_SIGNED(129,11),
TO_SIGNED(82,11),
TO_SIGNED(35,11),
TO_SIGNED(-12,11),
TO_SIGNED(-59,11),
TO_SIGNED(-105,11),
TO_SIGNED(-152,11),
TO_SIGNED(-197,11),
TO_SIGNED(-242,11),
TO_SIGNED(-286,11),
TO_SIGNED(-329,11),
TO_SIGNED(-371,11),
TO_SIGNED(-411,11),
TO_SIGNED(-449,11),
TO_SIGNED(-486,11),
TO_SIGNED(-521,11),
TO_SIGNED(-554,11),
TO_SIGNED(-584,11),
TO_SIGNED(-613,11),
TO_SIGNED(-639,11),
TO_SIGNED(-662,11),
TO_SIGNED(-683,11),
TO_SIGNED(-701,11),
TO_SIGNED(-716,11),
TO_SIGNED(-729,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-711,11),
TO_SIGNED(-694,11),
TO_SIGNED(-675,11),
TO_SIGNED(-653,11),
TO_SIGNED(-629,11),
TO_SIGNED(-602,11),
TO_SIGNED(-573,11),
TO_SIGNED(-541,11),
TO_SIGNED(-508,11),
TO_SIGNED(-472,11),
TO_SIGNED(-435,11),
TO_SIGNED(-396,11),
TO_SIGNED(-355,11),
TO_SIGNED(-313,11),
TO_SIGNED(-270,11),
TO_SIGNED(-225,11),
TO_SIGNED(-180,11),
TO_SIGNED(-134,11),
TO_SIGNED(-87,11),
TO_SIGNED(-41,11),
TO_SIGNED(6,11),
TO_SIGNED(53,11),
TO_SIGNED(100,11),
TO_SIGNED(147,11),
TO_SIGNED(192,11),
TO_SIGNED(237,11),
TO_SIGNED(281,11),
TO_SIGNED(324,11),
TO_SIGNED(366,11),
TO_SIGNED(406,11),
TO_SIGNED(445,11),
TO_SIGNED(482,11),
TO_SIGNED(517,11),
TO_SIGNED(550,11),
TO_SIGNED(581,11),
TO_SIGNED(610,11),
TO_SIGNED(636,11),
TO_SIGNED(659,11),
TO_SIGNED(681,11),
TO_SIGNED(699,11),
TO_SIGNED(715,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(712,11),
TO_SIGNED(696,11),
TO_SIGNED(677,11),
TO_SIGNED(656,11),
TO_SIGNED(632,11),
TO_SIGNED(605,11),
TO_SIGNED(576,11),
TO_SIGNED(545,11),
TO_SIGNED(512,11),
TO_SIGNED(476,11),
TO_SIGNED(439,11),
TO_SIGNED(400,11),
TO_SIGNED(360,11),
TO_SIGNED(318,11),
TO_SIGNED(275,11),
TO_SIGNED(230,11),
TO_SIGNED(185,11),
TO_SIGNED(139,11),
TO_SIGNED(93,11),
TO_SIGNED(46,11),
TO_SIGNED(-1,11),
TO_SIGNED(-48,11),
TO_SIGNED(-95,11),
TO_SIGNED(-141,11),
TO_SIGNED(-187,11),
TO_SIGNED(-232,11),
TO_SIGNED(-276,11),
TO_SIGNED(-320,11),
TO_SIGNED(-362,11),
TO_SIGNED(-402,11),
TO_SIGNED(-441,11),
TO_SIGNED(-478,11),
TO_SIGNED(-513,11),
TO_SIGNED(-547,11),
TO_SIGNED(-578,11),
TO_SIGNED(-606,11),
TO_SIGNED(-633,11),
TO_SIGNED(-657,11),
TO_SIGNED(-678,11),
TO_SIGNED(-697,11),
TO_SIGNED(-713,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-714,11),
TO_SIGNED(-698,11),
TO_SIGNED(-680,11),
TO_SIGNED(-658,11),
TO_SIGNED(-635,11),
TO_SIGNED(-608,11),
TO_SIGNED(-580,11),
TO_SIGNED(-549,11),
TO_SIGNED(-516,11),
TO_SIGNED(-480,11),
TO_SIGNED(-443,11),
TO_SIGNED(-405,11),
TO_SIGNED(-364,11),
TO_SIGNED(-323,11),
TO_SIGNED(-279,11),
TO_SIGNED(-235,11),
TO_SIGNED(-190,11),
TO_SIGNED(-144,11),
TO_SIGNED(-98,11),
TO_SIGNED(-51,11),
TO_SIGNED(-4,11),
TO_SIGNED(43,11),
TO_SIGNED(90,11),
TO_SIGNED(136,11),
TO_SIGNED(182,11),
TO_SIGNED(227,11),
TO_SIGNED(272,11),
TO_SIGNED(315,11),
TO_SIGNED(357,11),
TO_SIGNED(397,11),
TO_SIGNED(437,11),
TO_SIGNED(474,11),
TO_SIGNED(509,11),
TO_SIGNED(543,11),
TO_SIGNED(574,11),
TO_SIGNED(603,11),
TO_SIGNED(630,11),
TO_SIGNED(654,11),
TO_SIGNED(676,11),
TO_SIGNED(695,11),
TO_SIGNED(711,11),
TO_SIGNED(725,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(716,11),
TO_SIGNED(700,11),
TO_SIGNED(682,11),
TO_SIGNED(661,11),
TO_SIGNED(637,11),
TO_SIGNED(611,11),
TO_SIGNED(583,11),
TO_SIGNED(552,11),
TO_SIGNED(519,11),
TO_SIGNED(485,11),
TO_SIGNED(448,11),
TO_SIGNED(409,11),
TO_SIGNED(369,11),
TO_SIGNED(327,11),
TO_SIGNED(284,11),
TO_SIGNED(240,11),
TO_SIGNED(195,11),
TO_SIGNED(150,11),
TO_SIGNED(103,11),
TO_SIGNED(57,11),
TO_SIGNED(10,11),
TO_SIGNED(-37,11),
TO_SIGNED(-84,11),
TO_SIGNED(-131,11),
TO_SIGNED(-177,11),
TO_SIGNED(-222,11),
TO_SIGNED(-267,11),
TO_SIGNED(-310,11),
TO_SIGNED(-352,11),
TO_SIGNED(-393,11),
TO_SIGNED(-432,11),
TO_SIGNED(-470,11),
TO_SIGNED(-505,11),
TO_SIGNED(-539,11),
TO_SIGNED(-571,11),
TO_SIGNED(-600,11),
TO_SIGNED(-627,11),
TO_SIGNED(-652,11),
TO_SIGNED(-674,11),
TO_SIGNED(-693,11),
TO_SIGNED(-710,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-702,11),
TO_SIGNED(-684,11),
TO_SIGNED(-663,11),
TO_SIGNED(-640,11),
TO_SIGNED(-615,11),
TO_SIGNED(-586,11),
TO_SIGNED(-556,11),
TO_SIGNED(-523,11),
TO_SIGNED(-489,11),
TO_SIGNED(-452,11),
TO_SIGNED(-414,11),
TO_SIGNED(-374,11),
TO_SIGNED(-332,11),
TO_SIGNED(-289,11),
TO_SIGNED(-245,11),
TO_SIGNED(-201,11),
TO_SIGNED(-155,11),
TO_SIGNED(-109,11),
TO_SIGNED(-62,11),
TO_SIGNED(-15,11),
TO_SIGNED(32,11),
TO_SIGNED(79,11),
TO_SIGNED(125,11),
TO_SIGNED(172,11),
TO_SIGNED(217,11),
TO_SIGNED(262,11),
TO_SIGNED(305,11),
TO_SIGNED(347,11),
TO_SIGNED(388,11),
TO_SIGNED(428,11),
TO_SIGNED(466,11),
TO_SIGNED(501,11),
TO_SIGNED(535,11),
TO_SIGNED(567,11),
TO_SIGNED(597,11),
TO_SIGNED(624,11),
TO_SIGNED(649,11),
TO_SIGNED(671,11),
TO_SIGNED(691,11),
TO_SIGNED(708,11),
TO_SIGNED(722,11),
TO_SIGNED(733,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(704,11),
TO_SIGNED(686,11),
TO_SIGNED(666,11),
TO_SIGNED(643,11),
TO_SIGNED(618,11),
TO_SIGNED(590,11),
TO_SIGNED(559,11),
TO_SIGNED(527,11),
TO_SIGNED(493,11),
TO_SIGNED(456,11),
TO_SIGNED(418,11),
TO_SIGNED(378,11),
TO_SIGNED(337,11),
TO_SIGNED(294,11),
TO_SIGNED(250,11),
TO_SIGNED(206,11),
TO_SIGNED(160,11),
TO_SIGNED(114,11),
TO_SIGNED(67,11),
TO_SIGNED(20,11),
TO_SIGNED(-27,11),
TO_SIGNED(-74,11),
TO_SIGNED(-120,11),
TO_SIGNED(-166,11),
TO_SIGNED(-212,11),
TO_SIGNED(-257,11),
TO_SIGNED(-300,11),
TO_SIGNED(-343,11),
TO_SIGNED(-384,11),
TO_SIGNED(-423,11),
TO_SIGNED(-461,11),
TO_SIGNED(-497,11),
TO_SIGNED(-532,11),
TO_SIGNED(-564,11),
TO_SIGNED(-594,11),
TO_SIGNED(-621,11),
TO_SIGNED(-646,11),
TO_SIGNED(-669,11),
TO_SIGNED(-689,11),
TO_SIGNED(-706,11),
TO_SIGNED(-721,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-720,11),
TO_SIGNED(-706,11),
TO_SIGNED(-688,11),
TO_SIGNED(-668,11),
TO_SIGNED(-646,11),
TO_SIGNED(-621,11),
TO_SIGNED(-593,11),
TO_SIGNED(-563,11),
TO_SIGNED(-531,11),
TO_SIGNED(-497,11),
TO_SIGNED(-460,11),
TO_SIGNED(-422,11),
TO_SIGNED(-383,11),
TO_SIGNED(-342,11),
TO_SIGNED(-299,11),
TO_SIGNED(-256,11),
TO_SIGNED(-211,11),
TO_SIGNED(-165,11),
TO_SIGNED(-119,11),
TO_SIGNED(-73,11),
TO_SIGNED(-26,11),
TO_SIGNED(21,11),
TO_SIGNED(68,11),
TO_SIGNED(115,11),
TO_SIGNED(161,11),
TO_SIGNED(207,11),
TO_SIGNED(251,11),
TO_SIGNED(295,11),
TO_SIGNED(338,11),
TO_SIGNED(379,11),
TO_SIGNED(419,11),
TO_SIGNED(457,11),
TO_SIGNED(493,11),
TO_SIGNED(528,11),
TO_SIGNED(560,11),
TO_SIGNED(590,11),
TO_SIGNED(618,11),
TO_SIGNED(644,11),
TO_SIGNED(666,11),
TO_SIGNED(687,11),
TO_SIGNED(704,11),
TO_SIGNED(719,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(671,11),
TO_SIGNED(648,11),
TO_SIGNED(624,11),
TO_SIGNED(596,11),
TO_SIGNED(567,11),
TO_SIGNED(535,11),
TO_SIGNED(501,11),
TO_SIGNED(465,11),
TO_SIGNED(427,11),
TO_SIGNED(387,11),
TO_SIGNED(346,11),
TO_SIGNED(304,11),
TO_SIGNED(261,11),
TO_SIGNED(216,11),
TO_SIGNED(171,11),
TO_SIGNED(124,11),
TO_SIGNED(78,11),
TO_SIGNED(31,11),
TO_SIGNED(-16,11),
TO_SIGNED(-63,11),
TO_SIGNED(-110,11),
TO_SIGNED(-156,11),
TO_SIGNED(-202,11),
TO_SIGNED(-246,11),
TO_SIGNED(-290,11),
TO_SIGNED(-333,11),
TO_SIGNED(-375,11),
TO_SIGNED(-415,11),
TO_SIGNED(-453,11),
TO_SIGNED(-489,11),
TO_SIGNED(-524,11),
TO_SIGNED(-557,11),
TO_SIGNED(-587,11),
TO_SIGNED(-615,11),
TO_SIGNED(-641,11),
TO_SIGNED(-664,11),
TO_SIGNED(-685,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-730,11),
TO_SIGNED(-739,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-693,11),
TO_SIGNED(-673,11),
TO_SIGNED(-651,11),
TO_SIGNED(-627,11),
TO_SIGNED(-599,11),
TO_SIGNED(-570,11),
TO_SIGNED(-538,11),
TO_SIGNED(-505,11),
TO_SIGNED(-469,11),
TO_SIGNED(-431,11),
TO_SIGNED(-392,11),
TO_SIGNED(-351,11),
TO_SIGNED(-309,11),
TO_SIGNED(-266,11),
TO_SIGNED(-221,11),
TO_SIGNED(-176,11),
TO_SIGNED(-130,11),
TO_SIGNED(-83,11),
TO_SIGNED(-36,11),
TO_SIGNED(11,11),
TO_SIGNED(58,11),
TO_SIGNED(104,11),
TO_SIGNED(151,11),
TO_SIGNED(196,11),
TO_SIGNED(241,11),
TO_SIGNED(285,11),
TO_SIGNED(328,11),
TO_SIGNED(370,11),
TO_SIGNED(410,11),
TO_SIGNED(449,11),
TO_SIGNED(485,11),
TO_SIGNED(520,11),
TO_SIGNED(553,11),
TO_SIGNED(584,11),
TO_SIGNED(612,11),
TO_SIGNED(638,11),
TO_SIGNED(661,11),
TO_SIGNED(682,11),
TO_SIGNED(700,11),
TO_SIGNED(716,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(725,11),
TO_SIGNED(711,11),
TO_SIGNED(695,11),
TO_SIGNED(675,11),
TO_SIGNED(654,11),
TO_SIGNED(629,11),
TO_SIGNED(603,11),
TO_SIGNED(574,11),
TO_SIGNED(542,11),
TO_SIGNED(509,11),
TO_SIGNED(473,11),
TO_SIGNED(436,11),
TO_SIGNED(397,11),
TO_SIGNED(356,11),
TO_SIGNED(314,11),
TO_SIGNED(271,11),
TO_SIGNED(226,11),
TO_SIGNED(181,11),
TO_SIGNED(135,11),
TO_SIGNED(88,11),
TO_SIGNED(42,11),
TO_SIGNED(-5,11),
TO_SIGNED(-52,11),
TO_SIGNED(-99,11),
TO_SIGNED(-145,11),
TO_SIGNED(-191,11),
TO_SIGNED(-236,11),
TO_SIGNED(-280,11),
TO_SIGNED(-323,11),
TO_SIGNED(-365,11),
TO_SIGNED(-406,11),
TO_SIGNED(-444,11),
TO_SIGNED(-481,11),
TO_SIGNED(-516,11),
TO_SIGNED(-549,11),
TO_SIGNED(-580,11),
TO_SIGNED(-609,11),
TO_SIGNED(-635,11),
TO_SIGNED(-659,11),
TO_SIGNED(-680,11),
TO_SIGNED(-699,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-736,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-678,11),
TO_SIGNED(-656,11),
TO_SIGNED(-632,11),
TO_SIGNED(-606,11),
TO_SIGNED(-577,11),
TO_SIGNED(-546,11),
TO_SIGNED(-512,11),
TO_SIGNED(-477,11),
TO_SIGNED(-440,11),
TO_SIGNED(-401,11),
TO_SIGNED(-361,11),
TO_SIGNED(-319,11),
TO_SIGNED(-275,11),
TO_SIGNED(-231,11),
TO_SIGNED(-186,11),
TO_SIGNED(-140,11),
TO_SIGNED(-94,11),
TO_SIGNED(-47,11),
TO_SIGNED(0,11),
TO_SIGNED(47,11),
TO_SIGNED(94,11),
TO_SIGNED(140,11),
TO_SIGNED(186,11),
TO_SIGNED(231,11),
TO_SIGNED(275,11),
TO_SIGNED(319,11),
TO_SIGNED(361,11),
TO_SIGNED(401,11),
TO_SIGNED(440,11),
TO_SIGNED(477,11),
TO_SIGNED(512,11),
TO_SIGNED(546,11),
TO_SIGNED(577,11),
TO_SIGNED(606,11),
TO_SIGNED(632,11),
TO_SIGNED(656,11),
TO_SIGNED(678,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(736,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(699,11),
TO_SIGNED(680,11),
TO_SIGNED(659,11),
TO_SIGNED(635,11),
TO_SIGNED(609,11),
TO_SIGNED(580,11),
TO_SIGNED(549,11),
TO_SIGNED(516,11),
TO_SIGNED(481,11),
TO_SIGNED(444,11),
TO_SIGNED(406,11),
TO_SIGNED(365,11),
TO_SIGNED(323,11),
TO_SIGNED(280,11),
TO_SIGNED(236,11),
TO_SIGNED(191,11),
TO_SIGNED(145,11),
TO_SIGNED(99,11),
TO_SIGNED(52,11),
TO_SIGNED(5,11),
TO_SIGNED(-42,11),
TO_SIGNED(-88,11),
TO_SIGNED(-135,11),
TO_SIGNED(-181,11),
TO_SIGNED(-226,11),
TO_SIGNED(-271,11),
TO_SIGNED(-314,11),
TO_SIGNED(-356,11),
TO_SIGNED(-397,11),
TO_SIGNED(-436,11),
TO_SIGNED(-473,11),
TO_SIGNED(-509,11),
TO_SIGNED(-542,11),
TO_SIGNED(-574,11),
TO_SIGNED(-603,11),
TO_SIGNED(-629,11),
TO_SIGNED(-654,11),
TO_SIGNED(-675,11),
TO_SIGNED(-695,11),
TO_SIGNED(-711,11),
TO_SIGNED(-725,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-716,11),
TO_SIGNED(-700,11),
TO_SIGNED(-682,11),
TO_SIGNED(-661,11),
TO_SIGNED(-638,11),
TO_SIGNED(-612,11),
TO_SIGNED(-584,11),
TO_SIGNED(-553,11),
TO_SIGNED(-520,11),
TO_SIGNED(-485,11),
TO_SIGNED(-449,11),
TO_SIGNED(-410,11),
TO_SIGNED(-370,11),
TO_SIGNED(-328,11),
TO_SIGNED(-285,11),
TO_SIGNED(-241,11),
TO_SIGNED(-196,11),
TO_SIGNED(-151,11),
TO_SIGNED(-104,11),
TO_SIGNED(-58,11),
TO_SIGNED(-11,11),
TO_SIGNED(36,11),
TO_SIGNED(83,11),
TO_SIGNED(130,11),
TO_SIGNED(176,11),
TO_SIGNED(221,11),
TO_SIGNED(266,11),
TO_SIGNED(309,11),
TO_SIGNED(351,11),
TO_SIGNED(392,11),
TO_SIGNED(431,11),
TO_SIGNED(469,11),
TO_SIGNED(505,11),
TO_SIGNED(538,11),
TO_SIGNED(570,11),
TO_SIGNED(599,11),
TO_SIGNED(627,11),
TO_SIGNED(651,11),
TO_SIGNED(673,11),
TO_SIGNED(693,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(739,11),
TO_SIGNED(730,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(685,11),
TO_SIGNED(664,11),
TO_SIGNED(641,11),
TO_SIGNED(615,11),
TO_SIGNED(587,11),
TO_SIGNED(557,11),
TO_SIGNED(524,11),
TO_SIGNED(489,11),
TO_SIGNED(453,11),
TO_SIGNED(415,11),
TO_SIGNED(375,11),
TO_SIGNED(333,11),
TO_SIGNED(290,11),
TO_SIGNED(246,11),
TO_SIGNED(202,11),
TO_SIGNED(156,11),
TO_SIGNED(110,11),
TO_SIGNED(63,11),
TO_SIGNED(16,11),
TO_SIGNED(-31,11),
TO_SIGNED(-78,11),
TO_SIGNED(-124,11),
TO_SIGNED(-171,11),
TO_SIGNED(-216,11),
TO_SIGNED(-261,11),
TO_SIGNED(-304,11),
TO_SIGNED(-346,11),
TO_SIGNED(-387,11),
TO_SIGNED(-427,11),
TO_SIGNED(-465,11),
TO_SIGNED(-501,11),
TO_SIGNED(-535,11),
TO_SIGNED(-567,11),
TO_SIGNED(-596,11),
TO_SIGNED(-624,11),
TO_SIGNED(-648,11),
TO_SIGNED(-671,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-719,11),
TO_SIGNED(-704,11),
TO_SIGNED(-687,11),
TO_SIGNED(-666,11),
TO_SIGNED(-644,11),
TO_SIGNED(-618,11),
TO_SIGNED(-590,11),
TO_SIGNED(-560,11),
TO_SIGNED(-528,11),
TO_SIGNED(-493,11),
TO_SIGNED(-457,11),
TO_SIGNED(-419,11),
TO_SIGNED(-379,11),
TO_SIGNED(-338,11),
TO_SIGNED(-295,11),
TO_SIGNED(-251,11),
TO_SIGNED(-207,11),
TO_SIGNED(-161,11),
TO_SIGNED(-115,11),
TO_SIGNED(-68,11),
TO_SIGNED(-21,11),
TO_SIGNED(26,11),
TO_SIGNED(73,11),
TO_SIGNED(119,11),
TO_SIGNED(165,11),
TO_SIGNED(211,11),
TO_SIGNED(256,11),
TO_SIGNED(299,11),
TO_SIGNED(342,11),
TO_SIGNED(383,11),
TO_SIGNED(422,11),
TO_SIGNED(460,11),
TO_SIGNED(497,11),
TO_SIGNED(531,11),
TO_SIGNED(563,11),
TO_SIGNED(593,11),
TO_SIGNED(621,11),
TO_SIGNED(646,11),
TO_SIGNED(668,11),
TO_SIGNED(688,11),
TO_SIGNED(706,11),
TO_SIGNED(720,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(721,11),
TO_SIGNED(706,11),
TO_SIGNED(689,11),
TO_SIGNED(669,11),
TO_SIGNED(646,11),
TO_SIGNED(621,11),
TO_SIGNED(594,11),
TO_SIGNED(564,11),
TO_SIGNED(532,11),
TO_SIGNED(497,11),
TO_SIGNED(461,11),
TO_SIGNED(423,11),
TO_SIGNED(384,11),
TO_SIGNED(343,11),
TO_SIGNED(300,11),
TO_SIGNED(257,11),
TO_SIGNED(212,11),
TO_SIGNED(166,11),
TO_SIGNED(120,11),
TO_SIGNED(74,11),
TO_SIGNED(27,11),
TO_SIGNED(-20,11),
TO_SIGNED(-67,11),
TO_SIGNED(-114,11),
TO_SIGNED(-160,11),
TO_SIGNED(-206,11),
TO_SIGNED(-250,11),
TO_SIGNED(-294,11),
TO_SIGNED(-337,11),
TO_SIGNED(-378,11),
TO_SIGNED(-418,11),
TO_SIGNED(-456,11),
TO_SIGNED(-493,11),
TO_SIGNED(-527,11),
TO_SIGNED(-559,11),
TO_SIGNED(-590,11),
TO_SIGNED(-618,11),
TO_SIGNED(-643,11),
TO_SIGNED(-666,11),
TO_SIGNED(-686,11),
TO_SIGNED(-704,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-733,11),
TO_SIGNED(-722,11),
TO_SIGNED(-708,11),
TO_SIGNED(-691,11),
TO_SIGNED(-671,11),
TO_SIGNED(-649,11),
TO_SIGNED(-624,11),
TO_SIGNED(-597,11),
TO_SIGNED(-567,11),
TO_SIGNED(-535,11),
TO_SIGNED(-501,11),
TO_SIGNED(-466,11),
TO_SIGNED(-428,11),
TO_SIGNED(-388,11),
TO_SIGNED(-347,11),
TO_SIGNED(-305,11),
TO_SIGNED(-262,11),
TO_SIGNED(-217,11),
TO_SIGNED(-172,11),
TO_SIGNED(-125,11),
TO_SIGNED(-79,11),
TO_SIGNED(-32,11),
TO_SIGNED(15,11),
TO_SIGNED(62,11),
TO_SIGNED(109,11),
TO_SIGNED(155,11),
TO_SIGNED(201,11),
TO_SIGNED(245,11),
TO_SIGNED(289,11),
TO_SIGNED(332,11),
TO_SIGNED(374,11),
TO_SIGNED(414,11),
TO_SIGNED(452,11),
TO_SIGNED(489,11),
TO_SIGNED(523,11),
TO_SIGNED(556,11),
TO_SIGNED(586,11),
TO_SIGNED(615,11),
TO_SIGNED(640,11),
TO_SIGNED(663,11),
TO_SIGNED(684,11),
TO_SIGNED(702,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(710,11),
TO_SIGNED(693,11),
TO_SIGNED(674,11),
TO_SIGNED(652,11),
TO_SIGNED(627,11),
TO_SIGNED(600,11),
TO_SIGNED(571,11),
TO_SIGNED(539,11),
TO_SIGNED(505,11),
TO_SIGNED(470,11),
TO_SIGNED(432,11),
TO_SIGNED(393,11),
TO_SIGNED(352,11),
TO_SIGNED(310,11),
TO_SIGNED(267,11),
TO_SIGNED(222,11),
TO_SIGNED(177,11),
TO_SIGNED(131,11),
TO_SIGNED(84,11),
TO_SIGNED(37,11),
TO_SIGNED(-10,11),
TO_SIGNED(-57,11),
TO_SIGNED(-103,11),
TO_SIGNED(-150,11),
TO_SIGNED(-195,11),
TO_SIGNED(-240,11),
TO_SIGNED(-284,11),
TO_SIGNED(-327,11),
TO_SIGNED(-369,11),
TO_SIGNED(-409,11),
TO_SIGNED(-448,11),
TO_SIGNED(-485,11),
TO_SIGNED(-519,11),
TO_SIGNED(-552,11),
TO_SIGNED(-583,11),
TO_SIGNED(-611,11),
TO_SIGNED(-637,11),
TO_SIGNED(-661,11),
TO_SIGNED(-682,11),
TO_SIGNED(-700,11),
TO_SIGNED(-716,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-725,11),
TO_SIGNED(-711,11),
TO_SIGNED(-695,11),
TO_SIGNED(-676,11),
TO_SIGNED(-654,11),
TO_SIGNED(-630,11),
TO_SIGNED(-603,11),
TO_SIGNED(-574,11),
TO_SIGNED(-543,11),
TO_SIGNED(-509,11),
TO_SIGNED(-474,11),
TO_SIGNED(-437,11),
TO_SIGNED(-397,11),
TO_SIGNED(-357,11),
TO_SIGNED(-315,11),
TO_SIGNED(-272,11),
TO_SIGNED(-227,11),
TO_SIGNED(-182,11),
TO_SIGNED(-136,11),
TO_SIGNED(-90,11),
TO_SIGNED(-43,11),
TO_SIGNED(4,11),
TO_SIGNED(51,11),
TO_SIGNED(98,11),
TO_SIGNED(144,11),
TO_SIGNED(190,11),
TO_SIGNED(235,11),
TO_SIGNED(279,11),
TO_SIGNED(323,11),
TO_SIGNED(364,11),
TO_SIGNED(405,11),
TO_SIGNED(443,11),
TO_SIGNED(480,11),
TO_SIGNED(516,11),
TO_SIGNED(549,11),
TO_SIGNED(580,11),
TO_SIGNED(608,11),
TO_SIGNED(635,11),
TO_SIGNED(658,11),
TO_SIGNED(680,11),
TO_SIGNED(698,11),
TO_SIGNED(714,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(713,11),
TO_SIGNED(697,11),
TO_SIGNED(678,11),
TO_SIGNED(657,11),
TO_SIGNED(633,11),
TO_SIGNED(606,11),
TO_SIGNED(578,11),
TO_SIGNED(547,11),
TO_SIGNED(513,11),
TO_SIGNED(478,11),
TO_SIGNED(441,11),
TO_SIGNED(402,11),
TO_SIGNED(362,11),
TO_SIGNED(320,11),
TO_SIGNED(276,11),
TO_SIGNED(232,11),
TO_SIGNED(187,11),
TO_SIGNED(141,11),
TO_SIGNED(95,11),
TO_SIGNED(48,11),
TO_SIGNED(1,11),
TO_SIGNED(-46,11),
TO_SIGNED(-93,11),
TO_SIGNED(-139,11),
TO_SIGNED(-185,11),
TO_SIGNED(-230,11),
TO_SIGNED(-275,11),
TO_SIGNED(-318,11),
TO_SIGNED(-360,11),
TO_SIGNED(-400,11),
TO_SIGNED(-439,11),
TO_SIGNED(-476,11),
TO_SIGNED(-512,11),
TO_SIGNED(-545,11),
TO_SIGNED(-576,11),
TO_SIGNED(-605,11),
TO_SIGNED(-632,11),
TO_SIGNED(-656,11),
TO_SIGNED(-677,11),
TO_SIGNED(-696,11),
TO_SIGNED(-712,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-715,11),
TO_SIGNED(-699,11),
TO_SIGNED(-681,11),
TO_SIGNED(-659,11),
TO_SIGNED(-636,11),
TO_SIGNED(-610,11),
TO_SIGNED(-581,11),
TO_SIGNED(-550,11),
TO_SIGNED(-517,11),
TO_SIGNED(-482,11),
TO_SIGNED(-445,11),
TO_SIGNED(-406,11),
TO_SIGNED(-366,11),
TO_SIGNED(-324,11),
TO_SIGNED(-281,11),
TO_SIGNED(-237,11),
TO_SIGNED(-192,11),
TO_SIGNED(-147,11),
TO_SIGNED(-100,11),
TO_SIGNED(-53,11),
TO_SIGNED(-6,11),
TO_SIGNED(41,11),
TO_SIGNED(87,11),
TO_SIGNED(134,11),
TO_SIGNED(180,11),
TO_SIGNED(225,11),
TO_SIGNED(270,11),
TO_SIGNED(313,11),
TO_SIGNED(355,11),
TO_SIGNED(396,11),
TO_SIGNED(435,11),
TO_SIGNED(472,11),
TO_SIGNED(508,11),
TO_SIGNED(541,11),
TO_SIGNED(573,11),
TO_SIGNED(602,11),
TO_SIGNED(629,11),
TO_SIGNED(653,11),
TO_SIGNED(675,11),
TO_SIGNED(694,11),
TO_SIGNED(711,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(729,11),
TO_SIGNED(716,11),
TO_SIGNED(701,11),
TO_SIGNED(683,11),
TO_SIGNED(662,11),
TO_SIGNED(639,11),
TO_SIGNED(613,11),
TO_SIGNED(584,11),
TO_SIGNED(554,11),
TO_SIGNED(521,11),
TO_SIGNED(486,11),
TO_SIGNED(449,11),
TO_SIGNED(411,11),
TO_SIGNED(371,11),
TO_SIGNED(329,11),
TO_SIGNED(286,11),
TO_SIGNED(242,11),
TO_SIGNED(197,11),
TO_SIGNED(152,11),
TO_SIGNED(105,11),
TO_SIGNED(59,11),
TO_SIGNED(12,11),
TO_SIGNED(-35,11),
TO_SIGNED(-82,11),
TO_SIGNED(-129,11),
TO_SIGNED(-175,11),
TO_SIGNED(-220,11),
TO_SIGNED(-265,11),
TO_SIGNED(-308,11),
TO_SIGNED(-350,11),
TO_SIGNED(-391,11),
TO_SIGNED(-430,11),
TO_SIGNED(-468,11),
TO_SIGNED(-504,11),
TO_SIGNED(-538,11),
TO_SIGNED(-569,11),
TO_SIGNED(-599,11),
TO_SIGNED(-626,11),
TO_SIGNED(-651,11),
TO_SIGNED(-673,11),
TO_SIGNED(-692,11),
TO_SIGNED(-709,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-685,11),
TO_SIGNED(-664,11),
TO_SIGNED(-641,11),
TO_SIGNED(-616,11),
TO_SIGNED(-588,11),
TO_SIGNED(-557,11),
TO_SIGNED(-525,11),
TO_SIGNED(-490,11),
TO_SIGNED(-454,11),
TO_SIGNED(-415,11),
TO_SIGNED(-375,11),
TO_SIGNED(-334,11),
TO_SIGNED(-291,11),
TO_SIGNED(-247,11),
TO_SIGNED(-203,11),
TO_SIGNED(-157,11),
TO_SIGNED(-111,11),
TO_SIGNED(-64,11),
TO_SIGNED(-17,11),
TO_SIGNED(30,11),
TO_SIGNED(77,11),
TO_SIGNED(123,11),
TO_SIGNED(169,11),
TO_SIGNED(215,11),
TO_SIGNED(260,11),
TO_SIGNED(303,11),
TO_SIGNED(345,11),
TO_SIGNED(387,11),
TO_SIGNED(426,11),
TO_SIGNED(464,11),
TO_SIGNED(500,11),
TO_SIGNED(534,11),
TO_SIGNED(566,11),
TO_SIGNED(596,11),
TO_SIGNED(623,11),
TO_SIGNED(648,11),
TO_SIGNED(670,11),
TO_SIGNED(690,11),
TO_SIGNED(707,11),
TO_SIGNED(721,11),
TO_SIGNED(733,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(705,11),
TO_SIGNED(687,11),
TO_SIGNED(667,11),
TO_SIGNED(644,11),
TO_SIGNED(619,11),
TO_SIGNED(591,11),
TO_SIGNED(561,11),
TO_SIGNED(529,11),
TO_SIGNED(494,11),
TO_SIGNED(458,11),
TO_SIGNED(420,11),
TO_SIGNED(380,11),
TO_SIGNED(339,11),
TO_SIGNED(296,11),
TO_SIGNED(252,11),
TO_SIGNED(208,11),
TO_SIGNED(162,11),
TO_SIGNED(116,11),
TO_SIGNED(69,11),
TO_SIGNED(22,11),
TO_SIGNED(-25,11),
TO_SIGNED(-71,11),
TO_SIGNED(-118,11),
TO_SIGNED(-164,11),
TO_SIGNED(-210,11),
TO_SIGNED(-255,11),
TO_SIGNED(-298,11),
TO_SIGNED(-341,11),
TO_SIGNED(-382,11),
TO_SIGNED(-422,11),
TO_SIGNED(-460,11),
TO_SIGNED(-496,11),
TO_SIGNED(-530,11),
TO_SIGNED(-562,11),
TO_SIGNED(-592,11),
TO_SIGNED(-620,11),
TO_SIGNED(-645,11),
TO_SIGNED(-668,11),
TO_SIGNED(-688,11),
TO_SIGNED(-705,11),
TO_SIGNED(-720,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-721,11),
TO_SIGNED(-706,11),
TO_SIGNED(-689,11),
TO_SIGNED(-669,11),
TO_SIGNED(-647,11),
TO_SIGNED(-622,11),
TO_SIGNED(-594,11),
TO_SIGNED(-564,11),
TO_SIGNED(-532,11),
TO_SIGNED(-498,11),
TO_SIGNED(-462,11),
TO_SIGNED(-424,11),
TO_SIGNED(-385,11),
TO_SIGNED(-344,11),
TO_SIGNED(-301,11),
TO_SIGNED(-258,11),
TO_SIGNED(-213,11),
TO_SIGNED(-167,11),
TO_SIGNED(-121,11),
TO_SIGNED(-75,11),
TO_SIGNED(-28,11),
TO_SIGNED(19,11),
TO_SIGNED(66,11),
TO_SIGNED(113,11),
TO_SIGNED(159,11),
TO_SIGNED(205,11),
TO_SIGNED(249,11),
TO_SIGNED(293,11),
TO_SIGNED(336,11),
TO_SIGNED(377,11),
TO_SIGNED(417,11),
TO_SIGNED(455,11),
TO_SIGNED(492,11),
TO_SIGNED(526,11),
TO_SIGNED(559,11),
TO_SIGNED(589,11),
TO_SIGNED(617,11),
TO_SIGNED(642,11),
TO_SIGNED(665,11),
TO_SIGNED(686,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(708,11),
TO_SIGNED(691,11),
TO_SIGNED(672,11),
TO_SIGNED(650,11),
TO_SIGNED(625,11),
TO_SIGNED(598,11),
TO_SIGNED(568,11),
TO_SIGNED(536,11),
TO_SIGNED(502,11),
TO_SIGNED(466,11),
TO_SIGNED(429,11),
TO_SIGNED(389,11),
TO_SIGNED(348,11),
TO_SIGNED(306,11),
TO_SIGNED(263,11),
TO_SIGNED(218,11),
TO_SIGNED(173,11),
TO_SIGNED(127,11),
TO_SIGNED(80,11),
TO_SIGNED(33,11),
TO_SIGNED(-14,11),
TO_SIGNED(-61,11),
TO_SIGNED(-108,11),
TO_SIGNED(-154,11),
TO_SIGNED(-200,11),
TO_SIGNED(-244,11),
TO_SIGNED(-288,11),
TO_SIGNED(-331,11),
TO_SIGNED(-373,11),
TO_SIGNED(-413,11),
TO_SIGNED(-451,11),
TO_SIGNED(-488,11),
TO_SIGNED(-523,11),
TO_SIGNED(-555,11),
TO_SIGNED(-586,11),
TO_SIGNED(-614,11),
TO_SIGNED(-640,11),
TO_SIGNED(-663,11),
TO_SIGNED(-684,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-729,11),
TO_SIGNED(-739,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-710,11),
TO_SIGNED(-693,11),
TO_SIGNED(-674,11),
TO_SIGNED(-652,11),
TO_SIGNED(-628,11),
TO_SIGNED(-601,11),
TO_SIGNED(-571,11),
TO_SIGNED(-540,11),
TO_SIGNED(-506,11),
TO_SIGNED(-471,11),
TO_SIGNED(-433,11),
TO_SIGNED(-394,11),
TO_SIGNED(-353,11),
TO_SIGNED(-311,11),
TO_SIGNED(-268,11),
TO_SIGNED(-223,11),
TO_SIGNED(-178,11),
TO_SIGNED(-132,11),
TO_SIGNED(-85,11),
TO_SIGNED(-38,11),
TO_SIGNED(9,11),
TO_SIGNED(56,11),
TO_SIGNED(102,11),
TO_SIGNED(149,11),
TO_SIGNED(194,11),
TO_SIGNED(239,11),
TO_SIGNED(283,11),
TO_SIGNED(326,11),
TO_SIGNED(368,11),
TO_SIGNED(408,11),
TO_SIGNED(447,11),
TO_SIGNED(484,11),
TO_SIGNED(519,11),
TO_SIGNED(552,11),
TO_SIGNED(582,11),
TO_SIGNED(611,11),
TO_SIGNED(637,11),
TO_SIGNED(660,11),
TO_SIGNED(681,11),
TO_SIGNED(700,11),
TO_SIGNED(715,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(736,11),
TO_SIGNED(725,11),
TO_SIGNED(712,11),
TO_SIGNED(695,11),
TO_SIGNED(676,11),
TO_SIGNED(655,11),
TO_SIGNED(631,11),
TO_SIGNED(604,11),
TO_SIGNED(575,11),
TO_SIGNED(544,11),
TO_SIGNED(510,11),
TO_SIGNED(475,11),
TO_SIGNED(437,11),
TO_SIGNED(398,11),
TO_SIGNED(358,11),
TO_SIGNED(316,11),
TO_SIGNED(273,11),
TO_SIGNED(228,11),
TO_SIGNED(183,11),
TO_SIGNED(137,11),
TO_SIGNED(91,11),
TO_SIGNED(44,11),
TO_SIGNED(-3,11),
TO_SIGNED(-50,11),
TO_SIGNED(-97,11),
TO_SIGNED(-143,11),
TO_SIGNED(-189,11),
TO_SIGNED(-234,11),
TO_SIGNED(-278,11),
TO_SIGNED(-322,11),
TO_SIGNED(-363,11),
TO_SIGNED(-404,11),
TO_SIGNED(-443,11),
TO_SIGNED(-480,11),
TO_SIGNED(-515,11),
TO_SIGNED(-548,11),
TO_SIGNED(-579,11),
TO_SIGNED(-608,11),
TO_SIGNED(-634,11),
TO_SIGNED(-658,11),
TO_SIGNED(-679,11),
TO_SIGNED(-698,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-679,11),
TO_SIGNED(-657,11),
TO_SIGNED(-633,11),
TO_SIGNED(-607,11),
TO_SIGNED(-578,11),
TO_SIGNED(-547,11),
TO_SIGNED(-514,11),
TO_SIGNED(-479,11),
TO_SIGNED(-442,11),
TO_SIGNED(-403,11),
TO_SIGNED(-362,11),
TO_SIGNED(-321,11),
TO_SIGNED(-277,11),
TO_SIGNED(-233,11),
TO_SIGNED(-188,11),
TO_SIGNED(-142,11),
TO_SIGNED(-96,11),
TO_SIGNED(-49,11),
TO_SIGNED(-2,11),
TO_SIGNED(45,11),
TO_SIGNED(92,11),
TO_SIGNED(138,11),
TO_SIGNED(184,11),
TO_SIGNED(229,11),
TO_SIGNED(274,11),
TO_SIGNED(317,11),
TO_SIGNED(359,11),
TO_SIGNED(399,11),
TO_SIGNED(438,11),
TO_SIGNED(476,11),
TO_SIGNED(511,11),
TO_SIGNED(544,11),
TO_SIGNED(576,11),
TO_SIGNED(605,11),
TO_SIGNED(631,11),
TO_SIGNED(655,11),
TO_SIGNED(677,11),
TO_SIGNED(696,11),
TO_SIGNED(712,11),
TO_SIGNED(725,11),
TO_SIGNED(736,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(715,11),
TO_SIGNED(699,11),
TO_SIGNED(681,11),
TO_SIGNED(660,11),
TO_SIGNED(636,11),
TO_SIGNED(610,11),
TO_SIGNED(582,11),
TO_SIGNED(551,11),
TO_SIGNED(518,11),
TO_SIGNED(483,11),
TO_SIGNED(446,11),
TO_SIGNED(407,11),
TO_SIGNED(367,11),
TO_SIGNED(325,11),
TO_SIGNED(282,11),
TO_SIGNED(238,11),
TO_SIGNED(193,11),
TO_SIGNED(148,11),
TO_SIGNED(101,11),
TO_SIGNED(54,11),
TO_SIGNED(7,11),
TO_SIGNED(-40,11),
TO_SIGNED(-86,11),
TO_SIGNED(-133,11),
TO_SIGNED(-179,11),
TO_SIGNED(-224,11),
TO_SIGNED(-269,11),
TO_SIGNED(-312,11),
TO_SIGNED(-354,11),
TO_SIGNED(-395,11),
TO_SIGNED(-434,11),
TO_SIGNED(-471,11),
TO_SIGNED(-507,11),
TO_SIGNED(-541,11),
TO_SIGNED(-572,11),
TO_SIGNED(-601,11),
TO_SIGNED(-628,11),
TO_SIGNED(-653,11),
TO_SIGNED(-675,11),
TO_SIGNED(-694,11),
TO_SIGNED(-710,11),
TO_SIGNED(-724,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-701,11),
TO_SIGNED(-683,11),
TO_SIGNED(-662,11),
TO_SIGNED(-639,11),
TO_SIGNED(-613,11),
TO_SIGNED(-585,11),
TO_SIGNED(-554,11),
TO_SIGNED(-522,11),
TO_SIGNED(-487,11),
TO_SIGNED(-450,11),
TO_SIGNED(-412,11),
TO_SIGNED(-372,11),
TO_SIGNED(-330,11),
TO_SIGNED(-287,11),
TO_SIGNED(-243,11),
TO_SIGNED(-198,11),
TO_SIGNED(-153,11),
TO_SIGNED(-106,11),
TO_SIGNED(-60,11),
TO_SIGNED(-13,11),
TO_SIGNED(34,11),
TO_SIGNED(81,11),
TO_SIGNED(128,11),
TO_SIGNED(174,11),
TO_SIGNED(219,11),
TO_SIGNED(264,11),
TO_SIGNED(307,11),
TO_SIGNED(349,11),
TO_SIGNED(390,11),
TO_SIGNED(430,11),
TO_SIGNED(467,11),
TO_SIGNED(503,11),
TO_SIGNED(537,11),
TO_SIGNED(569,11),
TO_SIGNED(598,11),
TO_SIGNED(625,11),
TO_SIGNED(650,11),
TO_SIGNED(672,11),
TO_SIGNED(692,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(730,11),
TO_SIGNED(718,11),
TO_SIGNED(703,11),
TO_SIGNED(685,11),
TO_SIGNED(665,11),
TO_SIGNED(642,11),
TO_SIGNED(616,11),
TO_SIGNED(588,11),
TO_SIGNED(558,11),
TO_SIGNED(526,11),
TO_SIGNED(491,11),
TO_SIGNED(455,11),
TO_SIGNED(416,11),
TO_SIGNED(376,11),
TO_SIGNED(335,11),
TO_SIGNED(292,11),
TO_SIGNED(248,11),
TO_SIGNED(204,11),
TO_SIGNED(158,11),
TO_SIGNED(112,11),
TO_SIGNED(65,11),
TO_SIGNED(18,11),
TO_SIGNED(-29,11),
TO_SIGNED(-76,11),
TO_SIGNED(-122,11),
TO_SIGNED(-168,11),
TO_SIGNED(-214,11),
TO_SIGNED(-259,11),
TO_SIGNED(-302,11),
TO_SIGNED(-345,11),
TO_SIGNED(-386,11),
TO_SIGNED(-425,11),
TO_SIGNED(-463,11),
TO_SIGNED(-499,11),
TO_SIGNED(-533,11),
TO_SIGNED(-565,11),
TO_SIGNED(-595,11),
TO_SIGNED(-622,11),
TO_SIGNED(-647,11),
TO_SIGNED(-670,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-721,11),
TO_SIGNED(-733,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-720,11),
TO_SIGNED(-705,11),
TO_SIGNED(-688,11),
TO_SIGNED(-667,11),
TO_SIGNED(-645,11),
TO_SIGNED(-619,11),
TO_SIGNED(-592,11),
TO_SIGNED(-562,11),
TO_SIGNED(-529,11),
TO_SIGNED(-495,11),
TO_SIGNED(-459,11),
TO_SIGNED(-421,11),
TO_SIGNED(-381,11),
TO_SIGNED(-340,11),
TO_SIGNED(-297,11),
TO_SIGNED(-254,11),
TO_SIGNED(-209,11),
TO_SIGNED(-163,11),
TO_SIGNED(-117,11),
TO_SIGNED(-70,11),
TO_SIGNED(-24,11),
TO_SIGNED(24,11),
TO_SIGNED(70,11),
TO_SIGNED(117,11),
TO_SIGNED(163,11),
TO_SIGNED(209,11),
TO_SIGNED(254,11),
TO_SIGNED(297,11),
TO_SIGNED(340,11),
TO_SIGNED(381,11),
TO_SIGNED(421,11),
TO_SIGNED(459,11),
TO_SIGNED(495,11),
TO_SIGNED(529,11),
TO_SIGNED(562,11),
TO_SIGNED(592,11),
TO_SIGNED(619,11),
TO_SIGNED(645,11),
TO_SIGNED(667,11),
TO_SIGNED(688,11),
TO_SIGNED(705,11),
TO_SIGNED(720,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(733,11),
TO_SIGNED(721,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(670,11),
TO_SIGNED(647,11),
TO_SIGNED(622,11),
TO_SIGNED(595,11),
TO_SIGNED(565,11),
TO_SIGNED(533,11),
TO_SIGNED(499,11),
TO_SIGNED(463,11),
TO_SIGNED(425,11),
TO_SIGNED(386,11),
TO_SIGNED(345,11),
TO_SIGNED(302,11),
TO_SIGNED(259,11),
TO_SIGNED(214,11),
TO_SIGNED(168,11),
TO_SIGNED(122,11),
TO_SIGNED(76,11),
TO_SIGNED(29,11),
TO_SIGNED(-18,11),
TO_SIGNED(-65,11),
TO_SIGNED(-112,11),
TO_SIGNED(-158,11),
TO_SIGNED(-204,11),
TO_SIGNED(-248,11),
TO_SIGNED(-292,11),
TO_SIGNED(-335,11),
TO_SIGNED(-376,11),
TO_SIGNED(-416,11),
TO_SIGNED(-455,11),
TO_SIGNED(-491,11),
TO_SIGNED(-526,11),
TO_SIGNED(-558,11),
TO_SIGNED(-588,11),
TO_SIGNED(-616,11),
TO_SIGNED(-642,11),
TO_SIGNED(-665,11),
TO_SIGNED(-685,11),
TO_SIGNED(-703,11),
TO_SIGNED(-718,11),
TO_SIGNED(-730,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-692,11),
TO_SIGNED(-672,11),
TO_SIGNED(-650,11),
TO_SIGNED(-625,11),
TO_SIGNED(-598,11),
TO_SIGNED(-569,11),
TO_SIGNED(-537,11),
TO_SIGNED(-503,11),
TO_SIGNED(-467,11),
TO_SIGNED(-430,11),
TO_SIGNED(-390,11),
TO_SIGNED(-349,11),
TO_SIGNED(-307,11),
TO_SIGNED(-264,11),
TO_SIGNED(-219,11),
TO_SIGNED(-174,11),
TO_SIGNED(-128,11),
TO_SIGNED(-81,11),
TO_SIGNED(-34,11),
TO_SIGNED(13,11),
TO_SIGNED(60,11),
TO_SIGNED(106,11),
TO_SIGNED(153,11),
TO_SIGNED(198,11),
TO_SIGNED(243,11),
TO_SIGNED(287,11),
TO_SIGNED(330,11),
TO_SIGNED(372,11),
TO_SIGNED(412,11),
TO_SIGNED(450,11),
TO_SIGNED(487,11),
TO_SIGNED(522,11),
TO_SIGNED(554,11),
TO_SIGNED(585,11),
TO_SIGNED(613,11),
TO_SIGNED(639,11),
TO_SIGNED(662,11),
TO_SIGNED(683,11),
TO_SIGNED(701,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(724,11),
TO_SIGNED(710,11),
TO_SIGNED(694,11),
TO_SIGNED(675,11),
TO_SIGNED(653,11),
TO_SIGNED(628,11),
TO_SIGNED(601,11),
TO_SIGNED(572,11),
TO_SIGNED(541,11),
TO_SIGNED(507,11),
TO_SIGNED(471,11),
TO_SIGNED(434,11),
TO_SIGNED(395,11),
TO_SIGNED(354,11),
TO_SIGNED(312,11),
TO_SIGNED(269,11),
TO_SIGNED(224,11),
TO_SIGNED(179,11),
TO_SIGNED(133,11),
TO_SIGNED(86,11),
TO_SIGNED(40,11),
TO_SIGNED(-7,11),
TO_SIGNED(-54,11),
TO_SIGNED(-101,11),
TO_SIGNED(-148,11),
TO_SIGNED(-193,11),
TO_SIGNED(-238,11),
TO_SIGNED(-282,11),
TO_SIGNED(-325,11),
TO_SIGNED(-367,11),
TO_SIGNED(-407,11),
TO_SIGNED(-446,11),
TO_SIGNED(-483,11),
TO_SIGNED(-518,11),
TO_SIGNED(-551,11),
TO_SIGNED(-582,11),
TO_SIGNED(-610,11),
TO_SIGNED(-636,11),
TO_SIGNED(-660,11),
TO_SIGNED(-681,11),
TO_SIGNED(-699,11),
TO_SIGNED(-715,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-736,11),
TO_SIGNED(-725,11),
TO_SIGNED(-712,11),
TO_SIGNED(-696,11),
TO_SIGNED(-677,11),
TO_SIGNED(-655,11),
TO_SIGNED(-631,11),
TO_SIGNED(-605,11),
TO_SIGNED(-576,11),
TO_SIGNED(-544,11),
TO_SIGNED(-511,11),
TO_SIGNED(-476,11),
TO_SIGNED(-438,11),
TO_SIGNED(-399,11),
TO_SIGNED(-359,11),
TO_SIGNED(-317,11),
TO_SIGNED(-274,11),
TO_SIGNED(-229,11),
TO_SIGNED(-184,11),
TO_SIGNED(-138,11),
TO_SIGNED(-92,11),
TO_SIGNED(-45,11),
TO_SIGNED(2,11),
TO_SIGNED(49,11),
TO_SIGNED(96,11),
TO_SIGNED(142,11),
TO_SIGNED(188,11),
TO_SIGNED(233,11),
TO_SIGNED(277,11),
TO_SIGNED(321,11),
TO_SIGNED(362,11),
TO_SIGNED(403,11),
TO_SIGNED(442,11),
TO_SIGNED(479,11),
TO_SIGNED(514,11),
TO_SIGNED(547,11),
TO_SIGNED(578,11),
TO_SIGNED(607,11),
TO_SIGNED(633,11),
TO_SIGNED(657,11),
TO_SIGNED(679,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(698,11),
TO_SIGNED(679,11),
TO_SIGNED(658,11),
TO_SIGNED(634,11),
TO_SIGNED(608,11),
TO_SIGNED(579,11),
TO_SIGNED(548,11),
TO_SIGNED(515,11),
TO_SIGNED(480,11),
TO_SIGNED(443,11),
TO_SIGNED(404,11),
TO_SIGNED(363,11),
TO_SIGNED(322,11),
TO_SIGNED(278,11),
TO_SIGNED(234,11),
TO_SIGNED(189,11),
TO_SIGNED(143,11),
TO_SIGNED(97,11),
TO_SIGNED(50,11),
TO_SIGNED(3,11),
TO_SIGNED(-44,11),
TO_SIGNED(-91,11),
TO_SIGNED(-137,11),
TO_SIGNED(-183,11),
TO_SIGNED(-228,11),
TO_SIGNED(-273,11),
TO_SIGNED(-316,11),
TO_SIGNED(-358,11),
TO_SIGNED(-398,11),
TO_SIGNED(-437,11),
TO_SIGNED(-475,11),
TO_SIGNED(-510,11),
TO_SIGNED(-544,11),
TO_SIGNED(-575,11),
TO_SIGNED(-604,11),
TO_SIGNED(-631,11),
TO_SIGNED(-655,11),
TO_SIGNED(-676,11),
TO_SIGNED(-695,11),
TO_SIGNED(-712,11),
TO_SIGNED(-725,11),
TO_SIGNED(-736,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-715,11),
TO_SIGNED(-700,11),
TO_SIGNED(-681,11),
TO_SIGNED(-660,11),
TO_SIGNED(-637,11),
TO_SIGNED(-611,11),
TO_SIGNED(-582,11),
TO_SIGNED(-552,11),
TO_SIGNED(-519,11),
TO_SIGNED(-484,11),
TO_SIGNED(-447,11),
TO_SIGNED(-408,11),
TO_SIGNED(-368,11),
TO_SIGNED(-326,11),
TO_SIGNED(-283,11),
TO_SIGNED(-239,11),
TO_SIGNED(-194,11),
TO_SIGNED(-149,11),
TO_SIGNED(-102,11),
TO_SIGNED(-56,11),
TO_SIGNED(-9,11),
TO_SIGNED(38,11),
TO_SIGNED(85,11),
TO_SIGNED(132,11),
TO_SIGNED(178,11),
TO_SIGNED(223,11),
TO_SIGNED(268,11),
TO_SIGNED(311,11),
TO_SIGNED(353,11),
TO_SIGNED(394,11),
TO_SIGNED(433,11),
TO_SIGNED(471,11),
TO_SIGNED(506,11),
TO_SIGNED(540,11),
TO_SIGNED(571,11),
TO_SIGNED(601,11),
TO_SIGNED(628,11),
TO_SIGNED(652,11),
TO_SIGNED(674,11),
TO_SIGNED(693,11),
TO_SIGNED(710,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(739,11),
TO_SIGNED(729,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(684,11),
TO_SIGNED(663,11),
TO_SIGNED(640,11),
TO_SIGNED(614,11),
TO_SIGNED(586,11),
TO_SIGNED(555,11),
TO_SIGNED(523,11),
TO_SIGNED(488,11),
TO_SIGNED(451,11),
TO_SIGNED(413,11),
TO_SIGNED(373,11),
TO_SIGNED(331,11),
TO_SIGNED(288,11),
TO_SIGNED(244,11),
TO_SIGNED(200,11),
TO_SIGNED(154,11),
TO_SIGNED(108,11),
TO_SIGNED(61,11),
TO_SIGNED(14,11),
TO_SIGNED(-33,11),
TO_SIGNED(-80,11),
TO_SIGNED(-127,11),
TO_SIGNED(-173,11),
TO_SIGNED(-218,11),
TO_SIGNED(-263,11),
TO_SIGNED(-306,11),
TO_SIGNED(-348,11),
TO_SIGNED(-389,11),
TO_SIGNED(-429,11),
TO_SIGNED(-466,11),
TO_SIGNED(-502,11),
TO_SIGNED(-536,11),
TO_SIGNED(-568,11),
TO_SIGNED(-598,11),
TO_SIGNED(-625,11),
TO_SIGNED(-650,11),
TO_SIGNED(-672,11),
TO_SIGNED(-691,11),
TO_SIGNED(-708,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-686,11),
TO_SIGNED(-665,11),
TO_SIGNED(-642,11),
TO_SIGNED(-617,11),
TO_SIGNED(-589,11),
TO_SIGNED(-559,11),
TO_SIGNED(-526,11),
TO_SIGNED(-492,11),
TO_SIGNED(-455,11),
TO_SIGNED(-417,11),
TO_SIGNED(-377,11),
TO_SIGNED(-336,11),
TO_SIGNED(-293,11),
TO_SIGNED(-249,11),
TO_SIGNED(-205,11),
TO_SIGNED(-159,11),
TO_SIGNED(-113,11),
TO_SIGNED(-66,11),
TO_SIGNED(-19,11),
TO_SIGNED(28,11),
TO_SIGNED(75,11),
TO_SIGNED(121,11),
TO_SIGNED(167,11),
TO_SIGNED(213,11),
TO_SIGNED(258,11),
TO_SIGNED(301,11),
TO_SIGNED(344,11),
TO_SIGNED(385,11),
TO_SIGNED(424,11),
TO_SIGNED(462,11),
TO_SIGNED(498,11),
TO_SIGNED(532,11),
TO_SIGNED(564,11),
TO_SIGNED(594,11),
TO_SIGNED(622,11),
TO_SIGNED(647,11),
TO_SIGNED(669,11),
TO_SIGNED(689,11),
TO_SIGNED(706,11),
TO_SIGNED(721,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(720,11),
TO_SIGNED(705,11),
TO_SIGNED(688,11),
TO_SIGNED(668,11),
TO_SIGNED(645,11),
TO_SIGNED(620,11),
TO_SIGNED(592,11),
TO_SIGNED(562,11),
TO_SIGNED(530,11),
TO_SIGNED(496,11),
TO_SIGNED(460,11),
TO_SIGNED(422,11),
TO_SIGNED(382,11),
TO_SIGNED(341,11),
TO_SIGNED(298,11),
TO_SIGNED(255,11),
TO_SIGNED(210,11),
TO_SIGNED(164,11),
TO_SIGNED(118,11),
TO_SIGNED(71,11),
TO_SIGNED(25,11),
TO_SIGNED(-22,11),
TO_SIGNED(-69,11),
TO_SIGNED(-116,11),
TO_SIGNED(-162,11),
TO_SIGNED(-208,11),
TO_SIGNED(-252,11),
TO_SIGNED(-296,11),
TO_SIGNED(-339,11),
TO_SIGNED(-380,11),
TO_SIGNED(-420,11),
TO_SIGNED(-458,11),
TO_SIGNED(-494,11),
TO_SIGNED(-529,11),
TO_SIGNED(-561,11),
TO_SIGNED(-591,11),
TO_SIGNED(-619,11),
TO_SIGNED(-644,11),
TO_SIGNED(-667,11),
TO_SIGNED(-687,11),
TO_SIGNED(-705,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-733,11),
TO_SIGNED(-721,11),
TO_SIGNED(-707,11),
TO_SIGNED(-690,11),
TO_SIGNED(-670,11),
TO_SIGNED(-648,11),
TO_SIGNED(-623,11),
TO_SIGNED(-596,11),
TO_SIGNED(-566,11),
TO_SIGNED(-534,11),
TO_SIGNED(-500,11),
TO_SIGNED(-464,11),
TO_SIGNED(-426,11),
TO_SIGNED(-387,11),
TO_SIGNED(-345,11),
TO_SIGNED(-303,11),
TO_SIGNED(-260,11),
TO_SIGNED(-215,11),
TO_SIGNED(-169,11),
TO_SIGNED(-123,11),
TO_SIGNED(-77,11),
TO_SIGNED(-30,11),
TO_SIGNED(17,11),
TO_SIGNED(64,11),
TO_SIGNED(111,11),
TO_SIGNED(157,11),
TO_SIGNED(203,11),
TO_SIGNED(247,11),
TO_SIGNED(291,11),
TO_SIGNED(334,11),
TO_SIGNED(375,11),
TO_SIGNED(415,11),
TO_SIGNED(454,11),
TO_SIGNED(490,11),
TO_SIGNED(525,11),
TO_SIGNED(557,11),
TO_SIGNED(588,11),
TO_SIGNED(616,11),
TO_SIGNED(641,11),
TO_SIGNED(664,11),
TO_SIGNED(685,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(709,11),
TO_SIGNED(692,11),
TO_SIGNED(673,11),
TO_SIGNED(651,11),
TO_SIGNED(626,11),
TO_SIGNED(599,11),
TO_SIGNED(569,11),
TO_SIGNED(538,11),
TO_SIGNED(504,11),
TO_SIGNED(468,11),
TO_SIGNED(430,11),
TO_SIGNED(391,11),
TO_SIGNED(350,11),
TO_SIGNED(308,11),
TO_SIGNED(265,11),
TO_SIGNED(220,11),
TO_SIGNED(175,11),
TO_SIGNED(129,11),
TO_SIGNED(82,11),
TO_SIGNED(35,11),
TO_SIGNED(-12,11),
TO_SIGNED(-59,11),
TO_SIGNED(-105,11),
TO_SIGNED(-152,11),
TO_SIGNED(-197,11),
TO_SIGNED(-242,11),
TO_SIGNED(-286,11),
TO_SIGNED(-329,11),
TO_SIGNED(-371,11),
TO_SIGNED(-411,11),
TO_SIGNED(-449,11),
TO_SIGNED(-486,11),
TO_SIGNED(-521,11),
TO_SIGNED(-554,11),
TO_SIGNED(-584,11),
TO_SIGNED(-613,11),
TO_SIGNED(-639,11),
TO_SIGNED(-662,11),
TO_SIGNED(-683,11),
TO_SIGNED(-701,11),
TO_SIGNED(-716,11),
TO_SIGNED(-729,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-711,11),
TO_SIGNED(-694,11),
TO_SIGNED(-675,11),
TO_SIGNED(-653,11),
TO_SIGNED(-629,11),
TO_SIGNED(-602,11),
TO_SIGNED(-573,11),
TO_SIGNED(-541,11),
TO_SIGNED(-508,11),
TO_SIGNED(-472,11),
TO_SIGNED(-435,11),
TO_SIGNED(-396,11),
TO_SIGNED(-355,11),
TO_SIGNED(-313,11),
TO_SIGNED(-270,11),
TO_SIGNED(-225,11),
TO_SIGNED(-180,11),
TO_SIGNED(-134,11),
TO_SIGNED(-87,11),
TO_SIGNED(-41,11),
TO_SIGNED(6,11),
TO_SIGNED(53,11),
TO_SIGNED(100,11),
TO_SIGNED(147,11),
TO_SIGNED(192,11),
TO_SIGNED(237,11),
TO_SIGNED(281,11),
TO_SIGNED(324,11),
TO_SIGNED(366,11),
TO_SIGNED(406,11),
TO_SIGNED(445,11),
TO_SIGNED(482,11),
TO_SIGNED(517,11),
TO_SIGNED(550,11),
TO_SIGNED(581,11),
TO_SIGNED(610,11),
TO_SIGNED(636,11),
TO_SIGNED(659,11),
TO_SIGNED(681,11),
TO_SIGNED(699,11),
TO_SIGNED(715,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(712,11),
TO_SIGNED(696,11),
TO_SIGNED(677,11),
TO_SIGNED(656,11),
TO_SIGNED(632,11),
TO_SIGNED(605,11),
TO_SIGNED(576,11),
TO_SIGNED(545,11),
TO_SIGNED(512,11),
TO_SIGNED(476,11),
TO_SIGNED(439,11),
TO_SIGNED(400,11),
TO_SIGNED(360,11),
TO_SIGNED(318,11),
TO_SIGNED(275,11),
TO_SIGNED(230,11),
TO_SIGNED(185,11),
TO_SIGNED(139,11),
TO_SIGNED(93,11),
TO_SIGNED(46,11),
TO_SIGNED(-1,11),
TO_SIGNED(-48,11),
TO_SIGNED(-95,11),
TO_SIGNED(-141,11),
TO_SIGNED(-187,11),
TO_SIGNED(-232,11),
TO_SIGNED(-276,11),
TO_SIGNED(-320,11),
TO_SIGNED(-362,11),
TO_SIGNED(-402,11),
TO_SIGNED(-441,11),
TO_SIGNED(-478,11),
TO_SIGNED(-513,11),
TO_SIGNED(-547,11),
TO_SIGNED(-578,11),
TO_SIGNED(-606,11),
TO_SIGNED(-633,11),
TO_SIGNED(-657,11),
TO_SIGNED(-678,11),
TO_SIGNED(-697,11),
TO_SIGNED(-713,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-714,11),
TO_SIGNED(-698,11),
TO_SIGNED(-680,11),
TO_SIGNED(-658,11),
TO_SIGNED(-635,11),
TO_SIGNED(-608,11),
TO_SIGNED(-580,11),
TO_SIGNED(-549,11),
TO_SIGNED(-516,11),
TO_SIGNED(-480,11),
TO_SIGNED(-443,11),
TO_SIGNED(-405,11),
TO_SIGNED(-364,11),
TO_SIGNED(-323,11),
TO_SIGNED(-279,11),
TO_SIGNED(-235,11),
TO_SIGNED(-190,11),
TO_SIGNED(-144,11),
TO_SIGNED(-98,11),
TO_SIGNED(-51,11),
TO_SIGNED(-4,11),
TO_SIGNED(43,11),
TO_SIGNED(90,11),
TO_SIGNED(136,11),
TO_SIGNED(182,11),
TO_SIGNED(227,11),
TO_SIGNED(272,11),
TO_SIGNED(315,11),
TO_SIGNED(357,11),
TO_SIGNED(397,11),
TO_SIGNED(437,11),
TO_SIGNED(474,11),
TO_SIGNED(509,11),
TO_SIGNED(543,11),
TO_SIGNED(574,11),
TO_SIGNED(603,11),
TO_SIGNED(630,11),
TO_SIGNED(654,11),
TO_SIGNED(676,11),
TO_SIGNED(695,11),
TO_SIGNED(711,11),
TO_SIGNED(725,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(716,11),
TO_SIGNED(700,11),
TO_SIGNED(682,11),
TO_SIGNED(661,11),
TO_SIGNED(637,11),
TO_SIGNED(611,11),
TO_SIGNED(583,11),
TO_SIGNED(552,11),
TO_SIGNED(519,11),
TO_SIGNED(485,11),
TO_SIGNED(448,11),
TO_SIGNED(409,11),
TO_SIGNED(369,11),
TO_SIGNED(327,11),
TO_SIGNED(284,11),
TO_SIGNED(240,11),
TO_SIGNED(195,11),
TO_SIGNED(150,11),
TO_SIGNED(103,11),
TO_SIGNED(57,11),
TO_SIGNED(10,11),
TO_SIGNED(-37,11),
TO_SIGNED(-84,11),
TO_SIGNED(-131,11),
TO_SIGNED(-177,11),
TO_SIGNED(-222,11),
TO_SIGNED(-267,11),
TO_SIGNED(-310,11),
TO_SIGNED(-352,11),
TO_SIGNED(-393,11),
TO_SIGNED(-432,11),
TO_SIGNED(-470,11),
TO_SIGNED(-505,11),
TO_SIGNED(-539,11),
TO_SIGNED(-571,11),
TO_SIGNED(-600,11),
TO_SIGNED(-627,11),
TO_SIGNED(-652,11),
TO_SIGNED(-674,11),
TO_SIGNED(-693,11),
TO_SIGNED(-710,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-702,11),
TO_SIGNED(-684,11),
TO_SIGNED(-663,11),
TO_SIGNED(-640,11),
TO_SIGNED(-615,11),
TO_SIGNED(-586,11),
TO_SIGNED(-556,11),
TO_SIGNED(-523,11),
TO_SIGNED(-489,11),
TO_SIGNED(-452,11),
TO_SIGNED(-414,11),
TO_SIGNED(-374,11),
TO_SIGNED(-332,11),
TO_SIGNED(-289,11),
TO_SIGNED(-245,11),
TO_SIGNED(-201,11),
TO_SIGNED(-155,11),
TO_SIGNED(-109,11),
TO_SIGNED(-62,11),
TO_SIGNED(-15,11),
TO_SIGNED(32,11),
TO_SIGNED(79,11),
TO_SIGNED(125,11),
TO_SIGNED(172,11),
TO_SIGNED(217,11),
TO_SIGNED(262,11),
TO_SIGNED(305,11),
TO_SIGNED(347,11),
TO_SIGNED(388,11),
TO_SIGNED(428,11),
TO_SIGNED(466,11),
TO_SIGNED(501,11),
TO_SIGNED(535,11),
TO_SIGNED(567,11),
TO_SIGNED(597,11),
TO_SIGNED(624,11),
TO_SIGNED(649,11),
TO_SIGNED(671,11),
TO_SIGNED(691,11),
TO_SIGNED(708,11),
TO_SIGNED(722,11),
TO_SIGNED(733,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(704,11),
TO_SIGNED(686,11),
TO_SIGNED(666,11),
TO_SIGNED(643,11),
TO_SIGNED(618,11),
TO_SIGNED(590,11),
TO_SIGNED(559,11),
TO_SIGNED(527,11),
TO_SIGNED(493,11),
TO_SIGNED(456,11),
TO_SIGNED(418,11),
TO_SIGNED(378,11),
TO_SIGNED(337,11),
TO_SIGNED(294,11),
TO_SIGNED(250,11),
TO_SIGNED(206,11),
TO_SIGNED(160,11),
TO_SIGNED(114,11),
TO_SIGNED(67,11),
TO_SIGNED(20,11),
TO_SIGNED(-27,11),
TO_SIGNED(-74,11),
TO_SIGNED(-120,11),
TO_SIGNED(-166,11),
TO_SIGNED(-212,11),
TO_SIGNED(-257,11),
TO_SIGNED(-300,11),
TO_SIGNED(-343,11),
TO_SIGNED(-384,11),
TO_SIGNED(-423,11),
TO_SIGNED(-461,11),
TO_SIGNED(-497,11),
TO_SIGNED(-532,11),
TO_SIGNED(-564,11),
TO_SIGNED(-594,11),
TO_SIGNED(-621,11),
TO_SIGNED(-646,11),
TO_SIGNED(-669,11),
TO_SIGNED(-689,11),
TO_SIGNED(-706,11),
TO_SIGNED(-721,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-720,11),
TO_SIGNED(-706,11),
TO_SIGNED(-688,11),
TO_SIGNED(-668,11),
TO_SIGNED(-646,11),
TO_SIGNED(-621,11),
TO_SIGNED(-593,11),
TO_SIGNED(-563,11),
TO_SIGNED(-531,11),
TO_SIGNED(-497,11),
TO_SIGNED(-460,11),
TO_SIGNED(-422,11),
TO_SIGNED(-383,11),
TO_SIGNED(-342,11),
TO_SIGNED(-299,11),
TO_SIGNED(-256,11),
TO_SIGNED(-211,11),
TO_SIGNED(-165,11),
TO_SIGNED(-119,11),
TO_SIGNED(-73,11),
TO_SIGNED(-26,11),
TO_SIGNED(21,11),
TO_SIGNED(68,11),
TO_SIGNED(115,11),
TO_SIGNED(161,11),
TO_SIGNED(207,11),
TO_SIGNED(251,11),
TO_SIGNED(295,11),
TO_SIGNED(338,11),
TO_SIGNED(379,11),
TO_SIGNED(419,11),
TO_SIGNED(457,11),
TO_SIGNED(493,11),
TO_SIGNED(528,11),
TO_SIGNED(560,11),
TO_SIGNED(590,11),
TO_SIGNED(618,11),
TO_SIGNED(644,11),
TO_SIGNED(666,11),
TO_SIGNED(687,11),
TO_SIGNED(704,11),
TO_SIGNED(719,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(671,11),
TO_SIGNED(648,11),
TO_SIGNED(624,11),
TO_SIGNED(596,11),
TO_SIGNED(567,11),
TO_SIGNED(535,11),
TO_SIGNED(501,11),
TO_SIGNED(465,11),
TO_SIGNED(427,11),
TO_SIGNED(387,11),
TO_SIGNED(346,11),
TO_SIGNED(304,11),
TO_SIGNED(261,11),
TO_SIGNED(216,11),
TO_SIGNED(171,11),
TO_SIGNED(124,11),
TO_SIGNED(78,11),
TO_SIGNED(31,11),
TO_SIGNED(-16,11),
TO_SIGNED(-63,11),
TO_SIGNED(-110,11),
TO_SIGNED(-156,11),
TO_SIGNED(-202,11),
TO_SIGNED(-246,11),
TO_SIGNED(-290,11),
TO_SIGNED(-333,11),
TO_SIGNED(-375,11),
TO_SIGNED(-415,11),
TO_SIGNED(-453,11),
TO_SIGNED(-489,11),
TO_SIGNED(-524,11),
TO_SIGNED(-557,11),
TO_SIGNED(-587,11),
TO_SIGNED(-615,11),
TO_SIGNED(-641,11),
TO_SIGNED(-664,11),
TO_SIGNED(-685,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-730,11),
TO_SIGNED(-739,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-693,11),
TO_SIGNED(-673,11),
TO_SIGNED(-651,11),
TO_SIGNED(-627,11),
TO_SIGNED(-599,11),
TO_SIGNED(-570,11),
TO_SIGNED(-538,11),
TO_SIGNED(-505,11),
TO_SIGNED(-469,11),
TO_SIGNED(-431,11),
TO_SIGNED(-392,11),
TO_SIGNED(-351,11),
TO_SIGNED(-309,11),
TO_SIGNED(-266,11),
TO_SIGNED(-221,11),
TO_SIGNED(-176,11),
TO_SIGNED(-130,11),
TO_SIGNED(-83,11),
TO_SIGNED(-36,11),
TO_SIGNED(11,11),
TO_SIGNED(58,11),
TO_SIGNED(104,11),
TO_SIGNED(151,11),
TO_SIGNED(196,11),
TO_SIGNED(241,11),
TO_SIGNED(285,11),
TO_SIGNED(328,11),
TO_SIGNED(370,11),
TO_SIGNED(410,11),
TO_SIGNED(449,11),
TO_SIGNED(485,11),
TO_SIGNED(520,11),
TO_SIGNED(553,11),
TO_SIGNED(584,11),
TO_SIGNED(612,11),
TO_SIGNED(638,11),
TO_SIGNED(661,11),
TO_SIGNED(682,11),
TO_SIGNED(700,11),
TO_SIGNED(716,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(725,11),
TO_SIGNED(711,11),
TO_SIGNED(695,11),
TO_SIGNED(675,11),
TO_SIGNED(654,11),
TO_SIGNED(629,11),
TO_SIGNED(603,11),
TO_SIGNED(574,11),
TO_SIGNED(542,11),
TO_SIGNED(509,11),
TO_SIGNED(473,11),
TO_SIGNED(436,11),
TO_SIGNED(397,11),
TO_SIGNED(356,11),
TO_SIGNED(314,11),
TO_SIGNED(271,11),
TO_SIGNED(226,11),
TO_SIGNED(181,11),
TO_SIGNED(135,11),
TO_SIGNED(88,11),
TO_SIGNED(42,11),
TO_SIGNED(-5,11),
TO_SIGNED(-52,11),
TO_SIGNED(-99,11),
TO_SIGNED(-145,11),
TO_SIGNED(-191,11),
TO_SIGNED(-236,11),
TO_SIGNED(-280,11),
TO_SIGNED(-323,11),
TO_SIGNED(-365,11),
TO_SIGNED(-406,11),
TO_SIGNED(-444,11),
TO_SIGNED(-481,11),
TO_SIGNED(-516,11),
TO_SIGNED(-549,11),
TO_SIGNED(-580,11),
TO_SIGNED(-609,11),
TO_SIGNED(-635,11),
TO_SIGNED(-659,11),
TO_SIGNED(-680,11),
TO_SIGNED(-699,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-736,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-678,11),
TO_SIGNED(-656,11),
TO_SIGNED(-632,11),
TO_SIGNED(-606,11),
TO_SIGNED(-577,11),
TO_SIGNED(-546,11),
TO_SIGNED(-512,11),
TO_SIGNED(-477,11),
TO_SIGNED(-440,11),
TO_SIGNED(-401,11),
TO_SIGNED(-361,11),
TO_SIGNED(-319,11),
TO_SIGNED(-275,11),
TO_SIGNED(-231,11),
TO_SIGNED(-186,11),
TO_SIGNED(-140,11),
TO_SIGNED(-94,11),
TO_SIGNED(-47,11),
TO_SIGNED(0,11),
TO_SIGNED(47,11),
TO_SIGNED(94,11),
TO_SIGNED(140,11),
TO_SIGNED(186,11),
TO_SIGNED(231,11),
TO_SIGNED(275,11),
TO_SIGNED(319,11),
TO_SIGNED(361,11),
TO_SIGNED(401,11),
TO_SIGNED(440,11),
TO_SIGNED(477,11),
TO_SIGNED(512,11),
TO_SIGNED(546,11),
TO_SIGNED(577,11),
TO_SIGNED(606,11),
TO_SIGNED(632,11),
TO_SIGNED(656,11),
TO_SIGNED(678,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(736,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(699,11),
TO_SIGNED(680,11),
TO_SIGNED(659,11),
TO_SIGNED(635,11),
TO_SIGNED(609,11),
TO_SIGNED(580,11),
TO_SIGNED(549,11),
TO_SIGNED(516,11),
TO_SIGNED(481,11),
TO_SIGNED(444,11),
TO_SIGNED(406,11),
TO_SIGNED(365,11),
TO_SIGNED(323,11),
TO_SIGNED(280,11),
TO_SIGNED(236,11),
TO_SIGNED(191,11),
TO_SIGNED(145,11),
TO_SIGNED(99,11),
TO_SIGNED(52,11),
TO_SIGNED(5,11),
TO_SIGNED(-42,11),
TO_SIGNED(-88,11),
TO_SIGNED(-135,11),
TO_SIGNED(-181,11),
TO_SIGNED(-226,11),
TO_SIGNED(-271,11),
TO_SIGNED(-314,11),
TO_SIGNED(-356,11),
TO_SIGNED(-397,11),
TO_SIGNED(-436,11),
TO_SIGNED(-473,11),
TO_SIGNED(-509,11),
TO_SIGNED(-542,11),
TO_SIGNED(-574,11),
TO_SIGNED(-603,11),
TO_SIGNED(-629,11),
TO_SIGNED(-654,11),
TO_SIGNED(-675,11),
TO_SIGNED(-695,11),
TO_SIGNED(-711,11),
TO_SIGNED(-725,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-716,11),
TO_SIGNED(-700,11),
TO_SIGNED(-682,11),
TO_SIGNED(-661,11),
TO_SIGNED(-638,11),
TO_SIGNED(-612,11),
TO_SIGNED(-584,11),
TO_SIGNED(-553,11),
TO_SIGNED(-520,11),
TO_SIGNED(-485,11),
TO_SIGNED(-449,11),
TO_SIGNED(-410,11),
TO_SIGNED(-370,11),
TO_SIGNED(-328,11),
TO_SIGNED(-285,11),
TO_SIGNED(-241,11),
TO_SIGNED(-196,11),
TO_SIGNED(-151,11),
TO_SIGNED(-104,11),
TO_SIGNED(-58,11),
TO_SIGNED(-11,11),
TO_SIGNED(36,11),
TO_SIGNED(83,11),
TO_SIGNED(130,11),
TO_SIGNED(176,11),
TO_SIGNED(221,11),
TO_SIGNED(266,11),
TO_SIGNED(309,11),
TO_SIGNED(351,11),
TO_SIGNED(392,11),
TO_SIGNED(431,11),
TO_SIGNED(469,11),
TO_SIGNED(505,11),
TO_SIGNED(538,11),
TO_SIGNED(570,11),
TO_SIGNED(599,11),
TO_SIGNED(627,11),
TO_SIGNED(651,11),
TO_SIGNED(673,11),
TO_SIGNED(693,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(739,11),
TO_SIGNED(730,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(685,11),
TO_SIGNED(664,11),
TO_SIGNED(641,11),
TO_SIGNED(615,11),
TO_SIGNED(587,11),
TO_SIGNED(557,11),
TO_SIGNED(524,11),
TO_SIGNED(489,11),
TO_SIGNED(453,11),
TO_SIGNED(415,11),
TO_SIGNED(375,11),
TO_SIGNED(333,11),
TO_SIGNED(290,11),
TO_SIGNED(246,11),
TO_SIGNED(202,11),
TO_SIGNED(156,11),
TO_SIGNED(110,11),
TO_SIGNED(63,11),
TO_SIGNED(16,11),
TO_SIGNED(-31,11),
TO_SIGNED(-78,11),
TO_SIGNED(-124,11),
TO_SIGNED(-171,11),
TO_SIGNED(-216,11),
TO_SIGNED(-261,11),
TO_SIGNED(-304,11),
TO_SIGNED(-346,11),
TO_SIGNED(-387,11),
TO_SIGNED(-427,11),
TO_SIGNED(-465,11),
TO_SIGNED(-501,11),
TO_SIGNED(-535,11),
TO_SIGNED(-567,11),
TO_SIGNED(-596,11),
TO_SIGNED(-624,11),
TO_SIGNED(-648,11),
TO_SIGNED(-671,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-719,11),
TO_SIGNED(-704,11),
TO_SIGNED(-687,11),
TO_SIGNED(-666,11),
TO_SIGNED(-644,11),
TO_SIGNED(-618,11),
TO_SIGNED(-590,11),
TO_SIGNED(-560,11),
TO_SIGNED(-528,11),
TO_SIGNED(-493,11),
TO_SIGNED(-457,11),
TO_SIGNED(-419,11),
TO_SIGNED(-379,11),
TO_SIGNED(-338,11),
TO_SIGNED(-295,11),
TO_SIGNED(-251,11),
TO_SIGNED(-207,11),
TO_SIGNED(-161,11),
TO_SIGNED(-115,11),
TO_SIGNED(-68,11),
TO_SIGNED(-21,11),
TO_SIGNED(26,11),
TO_SIGNED(73,11),
TO_SIGNED(119,11),
TO_SIGNED(165,11),
TO_SIGNED(211,11),
TO_SIGNED(256,11),
TO_SIGNED(299,11),
TO_SIGNED(342,11),
TO_SIGNED(383,11),
TO_SIGNED(422,11),
TO_SIGNED(460,11),
TO_SIGNED(497,11),
TO_SIGNED(531,11),
TO_SIGNED(563,11),
TO_SIGNED(593,11),
TO_SIGNED(621,11),
TO_SIGNED(646,11),
TO_SIGNED(668,11),
TO_SIGNED(688,11),
TO_SIGNED(706,11),
TO_SIGNED(720,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(721,11),
TO_SIGNED(706,11),
TO_SIGNED(689,11),
TO_SIGNED(669,11),
TO_SIGNED(646,11),
TO_SIGNED(621,11),
TO_SIGNED(594,11),
TO_SIGNED(564,11),
TO_SIGNED(532,11),
TO_SIGNED(497,11),
TO_SIGNED(461,11),
TO_SIGNED(423,11),
TO_SIGNED(384,11),
TO_SIGNED(343,11),
TO_SIGNED(300,11),
TO_SIGNED(257,11),
TO_SIGNED(212,11),
TO_SIGNED(166,11),
TO_SIGNED(120,11),
TO_SIGNED(74,11),
TO_SIGNED(27,11),
TO_SIGNED(-20,11),
TO_SIGNED(-67,11),
TO_SIGNED(-114,11),
TO_SIGNED(-160,11),
TO_SIGNED(-206,11),
TO_SIGNED(-250,11),
TO_SIGNED(-294,11),
TO_SIGNED(-337,11),
TO_SIGNED(-378,11),
TO_SIGNED(-418,11),
TO_SIGNED(-456,11),
TO_SIGNED(-493,11),
TO_SIGNED(-527,11),
TO_SIGNED(-559,11),
TO_SIGNED(-590,11),
TO_SIGNED(-618,11),
TO_SIGNED(-643,11),
TO_SIGNED(-666,11),
TO_SIGNED(-686,11),
TO_SIGNED(-704,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-733,11),
TO_SIGNED(-722,11),
TO_SIGNED(-708,11),
TO_SIGNED(-691,11),
TO_SIGNED(-671,11),
TO_SIGNED(-649,11),
TO_SIGNED(-624,11),
TO_SIGNED(-597,11),
TO_SIGNED(-567,11),
TO_SIGNED(-535,11),
TO_SIGNED(-501,11),
TO_SIGNED(-466,11),
TO_SIGNED(-428,11),
TO_SIGNED(-388,11),
TO_SIGNED(-347,11),
TO_SIGNED(-305,11),
TO_SIGNED(-262,11),
TO_SIGNED(-217,11),
TO_SIGNED(-172,11),
TO_SIGNED(-125,11),
TO_SIGNED(-79,11),
TO_SIGNED(-32,11),
TO_SIGNED(15,11),
TO_SIGNED(62,11),
TO_SIGNED(109,11),
TO_SIGNED(155,11),
TO_SIGNED(201,11),
TO_SIGNED(245,11),
TO_SIGNED(289,11),
TO_SIGNED(332,11),
TO_SIGNED(374,11),
TO_SIGNED(414,11),
TO_SIGNED(452,11),
TO_SIGNED(489,11),
TO_SIGNED(523,11),
TO_SIGNED(556,11),
TO_SIGNED(586,11),
TO_SIGNED(615,11),
TO_SIGNED(640,11),
TO_SIGNED(663,11),
TO_SIGNED(684,11),
TO_SIGNED(702,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(710,11),
TO_SIGNED(693,11),
TO_SIGNED(674,11),
TO_SIGNED(652,11),
TO_SIGNED(627,11),
TO_SIGNED(600,11),
TO_SIGNED(571,11),
TO_SIGNED(539,11),
TO_SIGNED(505,11),
TO_SIGNED(470,11),
TO_SIGNED(432,11),
TO_SIGNED(393,11),
TO_SIGNED(352,11),
TO_SIGNED(310,11),
TO_SIGNED(267,11),
TO_SIGNED(222,11),
TO_SIGNED(177,11),
TO_SIGNED(131,11),
TO_SIGNED(84,11),
TO_SIGNED(37,11),
TO_SIGNED(-10,11),
TO_SIGNED(-57,11),
TO_SIGNED(-103,11),
TO_SIGNED(-150,11),
TO_SIGNED(-195,11),
TO_SIGNED(-240,11),
TO_SIGNED(-284,11),
TO_SIGNED(-327,11),
TO_SIGNED(-369,11),
TO_SIGNED(-409,11),
TO_SIGNED(-448,11),
TO_SIGNED(-485,11),
TO_SIGNED(-519,11),
TO_SIGNED(-552,11),
TO_SIGNED(-583,11),
TO_SIGNED(-611,11),
TO_SIGNED(-637,11),
TO_SIGNED(-661,11),
TO_SIGNED(-682,11),
TO_SIGNED(-700,11),
TO_SIGNED(-716,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-725,11),
TO_SIGNED(-711,11),
TO_SIGNED(-695,11),
TO_SIGNED(-676,11),
TO_SIGNED(-654,11),
TO_SIGNED(-630,11),
TO_SIGNED(-603,11),
TO_SIGNED(-574,11),
TO_SIGNED(-543,11),
TO_SIGNED(-509,11),
TO_SIGNED(-474,11),
TO_SIGNED(-437,11),
TO_SIGNED(-397,11),
TO_SIGNED(-357,11),
TO_SIGNED(-315,11),
TO_SIGNED(-272,11),
TO_SIGNED(-227,11),
TO_SIGNED(-182,11),
TO_SIGNED(-136,11),
TO_SIGNED(-90,11),
TO_SIGNED(-43,11),
TO_SIGNED(4,11),
TO_SIGNED(51,11),
TO_SIGNED(98,11),
TO_SIGNED(144,11),
TO_SIGNED(190,11),
TO_SIGNED(235,11),
TO_SIGNED(279,11),
TO_SIGNED(323,11),
TO_SIGNED(364,11),
TO_SIGNED(405,11),
TO_SIGNED(443,11),
TO_SIGNED(480,11),
TO_SIGNED(516,11),
TO_SIGNED(549,11),
TO_SIGNED(580,11),
TO_SIGNED(608,11),
TO_SIGNED(635,11),
TO_SIGNED(658,11),
TO_SIGNED(680,11),
TO_SIGNED(698,11),
TO_SIGNED(714,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(713,11),
TO_SIGNED(697,11),
TO_SIGNED(678,11),
TO_SIGNED(657,11),
TO_SIGNED(633,11),
TO_SIGNED(606,11),
TO_SIGNED(578,11),
TO_SIGNED(547,11),
TO_SIGNED(513,11),
TO_SIGNED(478,11),
TO_SIGNED(441,11),
TO_SIGNED(402,11),
TO_SIGNED(362,11),
TO_SIGNED(320,11),
TO_SIGNED(276,11),
TO_SIGNED(232,11),
TO_SIGNED(187,11),
TO_SIGNED(141,11),
TO_SIGNED(95,11),
TO_SIGNED(48,11),
TO_SIGNED(1,11),
TO_SIGNED(-46,11),
TO_SIGNED(-93,11),
TO_SIGNED(-139,11),
TO_SIGNED(-185,11),
TO_SIGNED(-230,11),
TO_SIGNED(-275,11),
TO_SIGNED(-318,11),
TO_SIGNED(-360,11),
TO_SIGNED(-400,11),
TO_SIGNED(-439,11),
TO_SIGNED(-476,11),
TO_SIGNED(-512,11),
TO_SIGNED(-545,11),
TO_SIGNED(-576,11),
TO_SIGNED(-605,11),
TO_SIGNED(-632,11),
TO_SIGNED(-656,11),
TO_SIGNED(-677,11),
TO_SIGNED(-696,11),
TO_SIGNED(-712,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-715,11),
TO_SIGNED(-699,11),
TO_SIGNED(-681,11),
TO_SIGNED(-659,11),
TO_SIGNED(-636,11),
TO_SIGNED(-610,11),
TO_SIGNED(-581,11),
TO_SIGNED(-550,11),
TO_SIGNED(-517,11),
TO_SIGNED(-482,11),
TO_SIGNED(-445,11),
TO_SIGNED(-406,11),
TO_SIGNED(-366,11),
TO_SIGNED(-324,11),
TO_SIGNED(-281,11),
TO_SIGNED(-237,11),
TO_SIGNED(-192,11),
TO_SIGNED(-147,11),
TO_SIGNED(-100,11),
TO_SIGNED(-53,11),
TO_SIGNED(-6,11),
TO_SIGNED(41,11),
TO_SIGNED(87,11),
TO_SIGNED(134,11),
TO_SIGNED(180,11),
TO_SIGNED(225,11),
TO_SIGNED(270,11),
TO_SIGNED(313,11),
TO_SIGNED(355,11),
TO_SIGNED(396,11),
TO_SIGNED(435,11),
TO_SIGNED(472,11),
TO_SIGNED(508,11),
TO_SIGNED(541,11),
TO_SIGNED(573,11),
TO_SIGNED(602,11),
TO_SIGNED(629,11),
TO_SIGNED(653,11),
TO_SIGNED(675,11),
TO_SIGNED(694,11),
TO_SIGNED(711,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(729,11),
TO_SIGNED(716,11),
TO_SIGNED(701,11),
TO_SIGNED(683,11),
TO_SIGNED(662,11),
TO_SIGNED(639,11),
TO_SIGNED(613,11),
TO_SIGNED(584,11),
TO_SIGNED(554,11),
TO_SIGNED(521,11),
TO_SIGNED(486,11),
TO_SIGNED(449,11),
TO_SIGNED(411,11),
TO_SIGNED(371,11),
TO_SIGNED(329,11),
TO_SIGNED(286,11),
TO_SIGNED(242,11),
TO_SIGNED(197,11),
TO_SIGNED(152,11),
TO_SIGNED(105,11),
TO_SIGNED(59,11),
TO_SIGNED(12,11),
TO_SIGNED(-35,11),
TO_SIGNED(-82,11),
TO_SIGNED(-129,11),
TO_SIGNED(-175,11),
TO_SIGNED(-220,11),
TO_SIGNED(-265,11),
TO_SIGNED(-308,11),
TO_SIGNED(-350,11),
TO_SIGNED(-391,11),
TO_SIGNED(-430,11),
TO_SIGNED(-468,11),
TO_SIGNED(-504,11),
TO_SIGNED(-538,11),
TO_SIGNED(-569,11),
TO_SIGNED(-599,11),
TO_SIGNED(-626,11),
TO_SIGNED(-651,11),
TO_SIGNED(-673,11),
TO_SIGNED(-692,11),
TO_SIGNED(-709,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-685,11),
TO_SIGNED(-664,11),
TO_SIGNED(-641,11),
TO_SIGNED(-616,11),
TO_SIGNED(-588,11),
TO_SIGNED(-557,11),
TO_SIGNED(-525,11),
TO_SIGNED(-490,11),
TO_SIGNED(-454,11),
TO_SIGNED(-415,11),
TO_SIGNED(-375,11),
TO_SIGNED(-334,11),
TO_SIGNED(-291,11),
TO_SIGNED(-247,11),
TO_SIGNED(-203,11),
TO_SIGNED(-157,11),
TO_SIGNED(-111,11),
TO_SIGNED(-64,11),
TO_SIGNED(-17,11),
TO_SIGNED(30,11),
TO_SIGNED(77,11),
TO_SIGNED(123,11),
TO_SIGNED(169,11),
TO_SIGNED(215,11),
TO_SIGNED(260,11),
TO_SIGNED(303,11),
TO_SIGNED(345,11),
TO_SIGNED(387,11),
TO_SIGNED(426,11),
TO_SIGNED(464,11),
TO_SIGNED(500,11),
TO_SIGNED(534,11),
TO_SIGNED(566,11),
TO_SIGNED(596,11),
TO_SIGNED(623,11),
TO_SIGNED(648,11),
TO_SIGNED(670,11),
TO_SIGNED(690,11),
TO_SIGNED(707,11),
TO_SIGNED(721,11),
TO_SIGNED(733,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(705,11),
TO_SIGNED(687,11),
TO_SIGNED(667,11),
TO_SIGNED(644,11),
TO_SIGNED(619,11),
TO_SIGNED(591,11),
TO_SIGNED(561,11),
TO_SIGNED(529,11),
TO_SIGNED(494,11),
TO_SIGNED(458,11),
TO_SIGNED(420,11),
TO_SIGNED(380,11),
TO_SIGNED(339,11),
TO_SIGNED(296,11),
TO_SIGNED(252,11),
TO_SIGNED(208,11),
TO_SIGNED(162,11),
TO_SIGNED(116,11),
TO_SIGNED(69,11),
TO_SIGNED(22,11),
TO_SIGNED(-25,11),
TO_SIGNED(-71,11),
TO_SIGNED(-118,11),
TO_SIGNED(-164,11),
TO_SIGNED(-210,11),
TO_SIGNED(-255,11),
TO_SIGNED(-298,11),
TO_SIGNED(-341,11),
TO_SIGNED(-382,11),
TO_SIGNED(-422,11),
TO_SIGNED(-460,11),
TO_SIGNED(-496,11),
TO_SIGNED(-530,11),
TO_SIGNED(-562,11),
TO_SIGNED(-592,11),
TO_SIGNED(-620,11),
TO_SIGNED(-645,11),
TO_SIGNED(-668,11),
TO_SIGNED(-688,11),
TO_SIGNED(-705,11),
TO_SIGNED(-720,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-721,11),
TO_SIGNED(-706,11),
TO_SIGNED(-689,11),
TO_SIGNED(-669,11),
TO_SIGNED(-647,11),
TO_SIGNED(-622,11),
TO_SIGNED(-594,11),
TO_SIGNED(-564,11),
TO_SIGNED(-532,11),
TO_SIGNED(-498,11),
TO_SIGNED(-462,11),
TO_SIGNED(-424,11),
TO_SIGNED(-385,11),
TO_SIGNED(-344,11),
TO_SIGNED(-301,11),
TO_SIGNED(-258,11),
TO_SIGNED(-213,11),
TO_SIGNED(-167,11),
TO_SIGNED(-121,11),
TO_SIGNED(-75,11),
TO_SIGNED(-28,11),
TO_SIGNED(19,11),
TO_SIGNED(66,11),
TO_SIGNED(113,11),
TO_SIGNED(159,11),
TO_SIGNED(205,11),
TO_SIGNED(249,11),
TO_SIGNED(293,11),
TO_SIGNED(336,11),
TO_SIGNED(377,11),
TO_SIGNED(417,11),
TO_SIGNED(455,11),
TO_SIGNED(492,11),
TO_SIGNED(526,11),
TO_SIGNED(559,11),
TO_SIGNED(589,11),
TO_SIGNED(617,11),
TO_SIGNED(642,11),
TO_SIGNED(665,11),
TO_SIGNED(686,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(708,11),
TO_SIGNED(691,11),
TO_SIGNED(672,11),
TO_SIGNED(650,11),
TO_SIGNED(625,11),
TO_SIGNED(598,11),
TO_SIGNED(568,11),
TO_SIGNED(536,11),
TO_SIGNED(502,11),
TO_SIGNED(466,11),
TO_SIGNED(429,11),
TO_SIGNED(389,11),
TO_SIGNED(348,11),
TO_SIGNED(306,11),
TO_SIGNED(263,11),
TO_SIGNED(218,11),
TO_SIGNED(173,11),
TO_SIGNED(127,11),
TO_SIGNED(80,11),
TO_SIGNED(33,11),
TO_SIGNED(-14,11),
TO_SIGNED(-61,11),
TO_SIGNED(-108,11),
TO_SIGNED(-154,11),
TO_SIGNED(-200,11),
TO_SIGNED(-244,11),
TO_SIGNED(-288,11),
TO_SIGNED(-331,11),
TO_SIGNED(-373,11),
TO_SIGNED(-413,11),
TO_SIGNED(-451,11),
TO_SIGNED(-488,11),
TO_SIGNED(-523,11),
TO_SIGNED(-555,11),
TO_SIGNED(-586,11),
TO_SIGNED(-614,11),
TO_SIGNED(-640,11),
TO_SIGNED(-663,11),
TO_SIGNED(-684,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-729,11),
TO_SIGNED(-739,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-710,11),
TO_SIGNED(-693,11),
TO_SIGNED(-674,11),
TO_SIGNED(-652,11),
TO_SIGNED(-628,11),
TO_SIGNED(-601,11),
TO_SIGNED(-571,11),
TO_SIGNED(-540,11),
TO_SIGNED(-506,11),
TO_SIGNED(-471,11),
TO_SIGNED(-433,11),
TO_SIGNED(-394,11),
TO_SIGNED(-353,11),
TO_SIGNED(-311,11),
TO_SIGNED(-268,11),
TO_SIGNED(-223,11),
TO_SIGNED(-178,11),
TO_SIGNED(-132,11),
TO_SIGNED(-85,11),
TO_SIGNED(-38,11),
TO_SIGNED(9,11),
TO_SIGNED(56,11),
TO_SIGNED(102,11),
TO_SIGNED(149,11),
TO_SIGNED(194,11),
TO_SIGNED(239,11),
TO_SIGNED(283,11),
TO_SIGNED(326,11),
TO_SIGNED(368,11),
TO_SIGNED(408,11),
TO_SIGNED(447,11),
TO_SIGNED(484,11),
TO_SIGNED(519,11),
TO_SIGNED(552,11),
TO_SIGNED(582,11),
TO_SIGNED(611,11),
TO_SIGNED(637,11),
TO_SIGNED(660,11),
TO_SIGNED(681,11),
TO_SIGNED(700,11),
TO_SIGNED(715,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(736,11),
TO_SIGNED(725,11),
TO_SIGNED(712,11),
TO_SIGNED(695,11),
TO_SIGNED(676,11),
TO_SIGNED(655,11),
TO_SIGNED(631,11),
TO_SIGNED(604,11),
TO_SIGNED(575,11),
TO_SIGNED(544,11),
TO_SIGNED(510,11),
TO_SIGNED(475,11),
TO_SIGNED(437,11),
TO_SIGNED(398,11),
TO_SIGNED(358,11),
TO_SIGNED(316,11),
TO_SIGNED(273,11),
TO_SIGNED(228,11),
TO_SIGNED(183,11),
TO_SIGNED(137,11),
TO_SIGNED(91,11),
TO_SIGNED(44,11),
TO_SIGNED(-3,11),
TO_SIGNED(-50,11),
TO_SIGNED(-97,11),
TO_SIGNED(-143,11),
TO_SIGNED(-189,11),
TO_SIGNED(-234,11),
TO_SIGNED(-278,11),
TO_SIGNED(-322,11),
TO_SIGNED(-363,11),
TO_SIGNED(-404,11),
TO_SIGNED(-443,11),
TO_SIGNED(-480,11),
TO_SIGNED(-515,11),
TO_SIGNED(-548,11),
TO_SIGNED(-579,11),
TO_SIGNED(-608,11),
TO_SIGNED(-634,11),
TO_SIGNED(-658,11),
TO_SIGNED(-679,11),
TO_SIGNED(-698,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-679,11),
TO_SIGNED(-657,11),
TO_SIGNED(-633,11),
TO_SIGNED(-607,11),
TO_SIGNED(-578,11),
TO_SIGNED(-547,11),
TO_SIGNED(-514,11),
TO_SIGNED(-479,11),
TO_SIGNED(-442,11),
TO_SIGNED(-403,11),
TO_SIGNED(-362,11),
TO_SIGNED(-321,11),
TO_SIGNED(-277,11),
TO_SIGNED(-233,11),
TO_SIGNED(-188,11),
TO_SIGNED(-142,11),
TO_SIGNED(-96,11),
TO_SIGNED(-49,11),
TO_SIGNED(-2,11),
TO_SIGNED(45,11),
TO_SIGNED(92,11),
TO_SIGNED(138,11),
TO_SIGNED(184,11),
TO_SIGNED(229,11),
TO_SIGNED(274,11),
TO_SIGNED(317,11),
TO_SIGNED(359,11),
TO_SIGNED(399,11),
TO_SIGNED(438,11),
TO_SIGNED(476,11),
TO_SIGNED(511,11),
TO_SIGNED(544,11),
TO_SIGNED(576,11),
TO_SIGNED(605,11),
TO_SIGNED(631,11),
TO_SIGNED(655,11),
TO_SIGNED(677,11),
TO_SIGNED(696,11),
TO_SIGNED(712,11),
TO_SIGNED(725,11),
TO_SIGNED(736,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(715,11),
TO_SIGNED(699,11),
TO_SIGNED(681,11),
TO_SIGNED(660,11),
TO_SIGNED(636,11),
TO_SIGNED(610,11),
TO_SIGNED(582,11),
TO_SIGNED(551,11),
TO_SIGNED(518,11),
TO_SIGNED(483,11),
TO_SIGNED(446,11),
TO_SIGNED(407,11),
TO_SIGNED(367,11),
TO_SIGNED(325,11),
TO_SIGNED(282,11),
TO_SIGNED(238,11),
TO_SIGNED(193,11),
TO_SIGNED(148,11),
TO_SIGNED(101,11),
TO_SIGNED(54,11),
TO_SIGNED(7,11),
TO_SIGNED(-40,11),
TO_SIGNED(-86,11),
TO_SIGNED(-133,11),
TO_SIGNED(-179,11),
TO_SIGNED(-224,11),
TO_SIGNED(-269,11),
TO_SIGNED(-312,11),
TO_SIGNED(-354,11),
TO_SIGNED(-395,11),
TO_SIGNED(-434,11),
TO_SIGNED(-471,11),
TO_SIGNED(-507,11),
TO_SIGNED(-541,11),
TO_SIGNED(-572,11),
TO_SIGNED(-601,11),
TO_SIGNED(-628,11),
TO_SIGNED(-653,11),
TO_SIGNED(-675,11),
TO_SIGNED(-694,11),
TO_SIGNED(-710,11),
TO_SIGNED(-724,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-701,11),
TO_SIGNED(-683,11),
TO_SIGNED(-662,11),
TO_SIGNED(-639,11),
TO_SIGNED(-613,11),
TO_SIGNED(-585,11),
TO_SIGNED(-554,11),
TO_SIGNED(-522,11),
TO_SIGNED(-487,11),
TO_SIGNED(-450,11),
TO_SIGNED(-412,11),
TO_SIGNED(-372,11),
TO_SIGNED(-330,11),
TO_SIGNED(-287,11),
TO_SIGNED(-243,11),
TO_SIGNED(-198,11),
TO_SIGNED(-153,11),
TO_SIGNED(-106,11),
TO_SIGNED(-60,11),
TO_SIGNED(-13,11),
TO_SIGNED(34,11),
TO_SIGNED(81,11),
TO_SIGNED(128,11),
TO_SIGNED(174,11),
TO_SIGNED(219,11),
TO_SIGNED(264,11),
TO_SIGNED(307,11),
TO_SIGNED(349,11),
TO_SIGNED(390,11),
TO_SIGNED(430,11),
TO_SIGNED(467,11),
TO_SIGNED(503,11),
TO_SIGNED(537,11),
TO_SIGNED(569,11),
TO_SIGNED(598,11),
TO_SIGNED(625,11),
TO_SIGNED(650,11),
TO_SIGNED(672,11),
TO_SIGNED(692,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(730,11),
TO_SIGNED(718,11),
TO_SIGNED(703,11),
TO_SIGNED(685,11),
TO_SIGNED(665,11),
TO_SIGNED(642,11),
TO_SIGNED(616,11),
TO_SIGNED(588,11),
TO_SIGNED(558,11),
TO_SIGNED(526,11),
TO_SIGNED(491,11),
TO_SIGNED(455,11),
TO_SIGNED(416,11),
TO_SIGNED(376,11),
TO_SIGNED(335,11),
TO_SIGNED(292,11),
TO_SIGNED(248,11),
TO_SIGNED(204,11),
TO_SIGNED(158,11),
TO_SIGNED(112,11),
TO_SIGNED(65,11),
TO_SIGNED(18,11),
TO_SIGNED(-29,11),
TO_SIGNED(-76,11),
TO_SIGNED(-122,11),
TO_SIGNED(-168,11),
TO_SIGNED(-214,11),
TO_SIGNED(-259,11),
TO_SIGNED(-302,11),
TO_SIGNED(-345,11),
TO_SIGNED(-386,11),
TO_SIGNED(-425,11),
TO_SIGNED(-463,11),
TO_SIGNED(-499,11),
TO_SIGNED(-533,11),
TO_SIGNED(-565,11),
TO_SIGNED(-595,11),
TO_SIGNED(-622,11),
TO_SIGNED(-647,11),
TO_SIGNED(-670,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-721,11),
TO_SIGNED(-733,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-720,11),
TO_SIGNED(-705,11),
TO_SIGNED(-688,11),
TO_SIGNED(-667,11),
TO_SIGNED(-645,11),
TO_SIGNED(-619,11),
TO_SIGNED(-592,11),
TO_SIGNED(-562,11),
TO_SIGNED(-529,11),
TO_SIGNED(-495,11),
TO_SIGNED(-459,11),
TO_SIGNED(-421,11),
TO_SIGNED(-381,11),
TO_SIGNED(-340,11),
TO_SIGNED(-297,11),
TO_SIGNED(-254,11),
TO_SIGNED(-209,11),
TO_SIGNED(-163,11),
TO_SIGNED(-117,11),
TO_SIGNED(-70,11),
TO_SIGNED(-24,11),
TO_SIGNED(24,11),
TO_SIGNED(70,11),
TO_SIGNED(117,11),
TO_SIGNED(163,11),
TO_SIGNED(209,11),
TO_SIGNED(254,11),
TO_SIGNED(297,11),
TO_SIGNED(340,11),
TO_SIGNED(381,11),
TO_SIGNED(421,11),
TO_SIGNED(459,11),
TO_SIGNED(495,11),
TO_SIGNED(529,11),
TO_SIGNED(562,11),
TO_SIGNED(592,11),
TO_SIGNED(619,11),
TO_SIGNED(645,11),
TO_SIGNED(667,11),
TO_SIGNED(688,11),
TO_SIGNED(705,11),
TO_SIGNED(720,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(733,11),
TO_SIGNED(721,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(670,11),
TO_SIGNED(647,11),
TO_SIGNED(622,11),
TO_SIGNED(595,11),
TO_SIGNED(565,11),
TO_SIGNED(533,11),
TO_SIGNED(499,11),
TO_SIGNED(463,11),
TO_SIGNED(425,11),
TO_SIGNED(386,11),
TO_SIGNED(345,11),
TO_SIGNED(302,11),
TO_SIGNED(259,11),
TO_SIGNED(214,11),
TO_SIGNED(168,11),
TO_SIGNED(122,11),
TO_SIGNED(76,11),
TO_SIGNED(29,11),
TO_SIGNED(-18,11),
TO_SIGNED(-65,11),
TO_SIGNED(-112,11),
TO_SIGNED(-158,11),
TO_SIGNED(-204,11),
TO_SIGNED(-248,11),
TO_SIGNED(-292,11),
TO_SIGNED(-335,11),
TO_SIGNED(-376,11),
TO_SIGNED(-416,11),
TO_SIGNED(-455,11),
TO_SIGNED(-491,11),
TO_SIGNED(-526,11),
TO_SIGNED(-558,11),
TO_SIGNED(-588,11),
TO_SIGNED(-616,11),
TO_SIGNED(-642,11),
TO_SIGNED(-665,11),
TO_SIGNED(-685,11),
TO_SIGNED(-703,11),
TO_SIGNED(-718,11),
TO_SIGNED(-730,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-692,11),
TO_SIGNED(-672,11),
TO_SIGNED(-650,11),
TO_SIGNED(-625,11),
TO_SIGNED(-598,11),
TO_SIGNED(-569,11),
TO_SIGNED(-537,11),
TO_SIGNED(-503,11),
TO_SIGNED(-467,11),
TO_SIGNED(-430,11),
TO_SIGNED(-390,11),
TO_SIGNED(-349,11),
TO_SIGNED(-307,11),
TO_SIGNED(-264,11),
TO_SIGNED(-219,11),
TO_SIGNED(-174,11),
TO_SIGNED(-128,11),
TO_SIGNED(-81,11),
TO_SIGNED(-34,11),
TO_SIGNED(13,11),
TO_SIGNED(60,11),
TO_SIGNED(106,11),
TO_SIGNED(153,11),
TO_SIGNED(198,11),
TO_SIGNED(243,11),
TO_SIGNED(287,11),
TO_SIGNED(330,11),
TO_SIGNED(372,11),
TO_SIGNED(412,11),
TO_SIGNED(450,11),
TO_SIGNED(487,11),
TO_SIGNED(522,11),
TO_SIGNED(554,11),
TO_SIGNED(585,11),
TO_SIGNED(613,11),
TO_SIGNED(639,11),
TO_SIGNED(662,11),
TO_SIGNED(683,11),
TO_SIGNED(701,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(724,11),
TO_SIGNED(710,11),
TO_SIGNED(694,11),
TO_SIGNED(675,11),
TO_SIGNED(653,11),
TO_SIGNED(628,11),
TO_SIGNED(601,11),
TO_SIGNED(572,11),
TO_SIGNED(541,11),
TO_SIGNED(507,11),
TO_SIGNED(471,11),
TO_SIGNED(434,11),
TO_SIGNED(395,11),
TO_SIGNED(354,11),
TO_SIGNED(312,11),
TO_SIGNED(269,11),
TO_SIGNED(224,11),
TO_SIGNED(179,11),
TO_SIGNED(133,11),
TO_SIGNED(86,11),
TO_SIGNED(40,11),
TO_SIGNED(-7,11),
TO_SIGNED(-54,11),
TO_SIGNED(-101,11),
TO_SIGNED(-148,11),
TO_SIGNED(-193,11),
TO_SIGNED(-238,11),
TO_SIGNED(-282,11),
TO_SIGNED(-325,11),
TO_SIGNED(-367,11),
TO_SIGNED(-407,11),
TO_SIGNED(-446,11),
TO_SIGNED(-483,11),
TO_SIGNED(-518,11),
TO_SIGNED(-551,11),
TO_SIGNED(-582,11),
TO_SIGNED(-610,11),
TO_SIGNED(-636,11),
TO_SIGNED(-660,11),
TO_SIGNED(-681,11),
TO_SIGNED(-699,11),
TO_SIGNED(-715,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-736,11),
TO_SIGNED(-725,11),
TO_SIGNED(-712,11),
TO_SIGNED(-696,11),
TO_SIGNED(-677,11),
TO_SIGNED(-655,11),
TO_SIGNED(-631,11),
TO_SIGNED(-605,11),
TO_SIGNED(-576,11),
TO_SIGNED(-544,11),
TO_SIGNED(-511,11),
TO_SIGNED(-476,11),
TO_SIGNED(-438,11),
TO_SIGNED(-399,11),
TO_SIGNED(-359,11),
TO_SIGNED(-317,11),
TO_SIGNED(-274,11),
TO_SIGNED(-229,11),
TO_SIGNED(-184,11),
TO_SIGNED(-138,11),
TO_SIGNED(-92,11),
TO_SIGNED(-45,11),
TO_SIGNED(2,11),
TO_SIGNED(49,11),
TO_SIGNED(96,11),
TO_SIGNED(142,11),
TO_SIGNED(188,11),
TO_SIGNED(233,11),
TO_SIGNED(277,11),
TO_SIGNED(321,11),
TO_SIGNED(362,11),
TO_SIGNED(403,11),
TO_SIGNED(442,11),
TO_SIGNED(479,11),
TO_SIGNED(514,11),
TO_SIGNED(547,11),
TO_SIGNED(578,11),
TO_SIGNED(607,11),
TO_SIGNED(633,11),
TO_SIGNED(657,11),
TO_SIGNED(679,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(698,11),
TO_SIGNED(679,11),
TO_SIGNED(658,11),
TO_SIGNED(634,11),
TO_SIGNED(608,11),
TO_SIGNED(579,11),
TO_SIGNED(548,11),
TO_SIGNED(515,11),
TO_SIGNED(480,11),
TO_SIGNED(443,11),
TO_SIGNED(404,11),
TO_SIGNED(363,11),
TO_SIGNED(322,11),
TO_SIGNED(278,11),
TO_SIGNED(234,11),
TO_SIGNED(189,11),
TO_SIGNED(143,11),
TO_SIGNED(97,11),
TO_SIGNED(50,11),
TO_SIGNED(3,11),
TO_SIGNED(-44,11),
TO_SIGNED(-91,11),
TO_SIGNED(-137,11),
TO_SIGNED(-183,11),
TO_SIGNED(-228,11),
TO_SIGNED(-273,11),
TO_SIGNED(-316,11),
TO_SIGNED(-358,11),
TO_SIGNED(-398,11),
TO_SIGNED(-437,11),
TO_SIGNED(-475,11),
TO_SIGNED(-510,11),
TO_SIGNED(-544,11),
TO_SIGNED(-575,11),
TO_SIGNED(-604,11),
TO_SIGNED(-631,11),
TO_SIGNED(-655,11),
TO_SIGNED(-676,11),
TO_SIGNED(-695,11),
TO_SIGNED(-712,11),
TO_SIGNED(-725,11),
TO_SIGNED(-736,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-715,11),
TO_SIGNED(-700,11),
TO_SIGNED(-681,11),
TO_SIGNED(-660,11),
TO_SIGNED(-637,11),
TO_SIGNED(-611,11),
TO_SIGNED(-582,11),
TO_SIGNED(-552,11),
TO_SIGNED(-519,11),
TO_SIGNED(-484,11),
TO_SIGNED(-447,11),
TO_SIGNED(-408,11),
TO_SIGNED(-368,11),
TO_SIGNED(-326,11),
TO_SIGNED(-283,11),
TO_SIGNED(-239,11),
TO_SIGNED(-194,11),
TO_SIGNED(-149,11),
TO_SIGNED(-102,11),
TO_SIGNED(-56,11),
TO_SIGNED(-9,11),
TO_SIGNED(38,11),
TO_SIGNED(85,11),
TO_SIGNED(132,11),
TO_SIGNED(178,11),
TO_SIGNED(223,11),
TO_SIGNED(268,11),
TO_SIGNED(311,11),
TO_SIGNED(353,11),
TO_SIGNED(394,11),
TO_SIGNED(433,11),
TO_SIGNED(471,11),
TO_SIGNED(506,11),
TO_SIGNED(540,11),
TO_SIGNED(571,11),
TO_SIGNED(601,11),
TO_SIGNED(628,11),
TO_SIGNED(652,11),
TO_SIGNED(674,11),
TO_SIGNED(693,11),
TO_SIGNED(710,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(739,11),
TO_SIGNED(729,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(684,11),
TO_SIGNED(663,11),
TO_SIGNED(640,11),
TO_SIGNED(614,11),
TO_SIGNED(586,11),
TO_SIGNED(555,11),
TO_SIGNED(523,11),
TO_SIGNED(488,11),
TO_SIGNED(451,11),
TO_SIGNED(413,11),
TO_SIGNED(373,11),
TO_SIGNED(331,11),
TO_SIGNED(288,11),
TO_SIGNED(244,11),
TO_SIGNED(200,11),
TO_SIGNED(154,11),
TO_SIGNED(108,11),
TO_SIGNED(61,11),
TO_SIGNED(14,11),
TO_SIGNED(-33,11),
TO_SIGNED(-80,11),
TO_SIGNED(-127,11),
TO_SIGNED(-173,11),
TO_SIGNED(-218,11),
TO_SIGNED(-263,11),
TO_SIGNED(-306,11),
TO_SIGNED(-348,11),
TO_SIGNED(-389,11),
TO_SIGNED(-429,11),
TO_SIGNED(-466,11),
TO_SIGNED(-502,11),
TO_SIGNED(-536,11),
TO_SIGNED(-568,11),
TO_SIGNED(-598,11),
TO_SIGNED(-625,11),
TO_SIGNED(-650,11),
TO_SIGNED(-672,11),
TO_SIGNED(-691,11),
TO_SIGNED(-708,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-686,11),
TO_SIGNED(-665,11),
TO_SIGNED(-642,11),
TO_SIGNED(-617,11),
TO_SIGNED(-589,11),
TO_SIGNED(-559,11),
TO_SIGNED(-526,11),
TO_SIGNED(-492,11),
TO_SIGNED(-455,11),
TO_SIGNED(-417,11),
TO_SIGNED(-377,11),
TO_SIGNED(-336,11),
TO_SIGNED(-293,11),
TO_SIGNED(-249,11),
TO_SIGNED(-205,11),
TO_SIGNED(-159,11),
TO_SIGNED(-113,11),
TO_SIGNED(-66,11),
TO_SIGNED(-19,11),
TO_SIGNED(28,11),
TO_SIGNED(75,11),
TO_SIGNED(121,11),
TO_SIGNED(167,11),
TO_SIGNED(213,11),
TO_SIGNED(258,11),
TO_SIGNED(301,11),
TO_SIGNED(344,11),
TO_SIGNED(385,11),
TO_SIGNED(424,11),
TO_SIGNED(462,11),
TO_SIGNED(498,11),
TO_SIGNED(532,11),
TO_SIGNED(564,11),
TO_SIGNED(594,11),
TO_SIGNED(622,11),
TO_SIGNED(647,11),
TO_SIGNED(669,11),
TO_SIGNED(689,11),
TO_SIGNED(706,11),
TO_SIGNED(721,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(720,11),
TO_SIGNED(705,11),
TO_SIGNED(688,11),
TO_SIGNED(668,11),
TO_SIGNED(645,11),
TO_SIGNED(620,11),
TO_SIGNED(592,11),
TO_SIGNED(562,11),
TO_SIGNED(530,11),
TO_SIGNED(496,11),
TO_SIGNED(460,11),
TO_SIGNED(422,11),
TO_SIGNED(382,11),
TO_SIGNED(341,11),
TO_SIGNED(298,11),
TO_SIGNED(255,11),
TO_SIGNED(210,11),
TO_SIGNED(164,11),
TO_SIGNED(118,11),
TO_SIGNED(71,11),
TO_SIGNED(25,11),
TO_SIGNED(-22,11),
TO_SIGNED(-69,11),
TO_SIGNED(-116,11),
TO_SIGNED(-162,11),
TO_SIGNED(-208,11),
TO_SIGNED(-252,11),
TO_SIGNED(-296,11),
TO_SIGNED(-339,11),
TO_SIGNED(-380,11),
TO_SIGNED(-420,11),
TO_SIGNED(-458,11),
TO_SIGNED(-494,11),
TO_SIGNED(-529,11),
TO_SIGNED(-561,11),
TO_SIGNED(-591,11),
TO_SIGNED(-619,11),
TO_SIGNED(-644,11),
TO_SIGNED(-667,11),
TO_SIGNED(-687,11),
TO_SIGNED(-705,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-733,11),
TO_SIGNED(-721,11),
TO_SIGNED(-707,11),
TO_SIGNED(-690,11),
TO_SIGNED(-670,11),
TO_SIGNED(-648,11),
TO_SIGNED(-623,11),
TO_SIGNED(-596,11),
TO_SIGNED(-566,11),
TO_SIGNED(-534,11),
TO_SIGNED(-500,11),
TO_SIGNED(-464,11),
TO_SIGNED(-426,11),
TO_SIGNED(-387,11),
TO_SIGNED(-345,11),
TO_SIGNED(-303,11),
TO_SIGNED(-260,11),
TO_SIGNED(-215,11),
TO_SIGNED(-169,11),
TO_SIGNED(-123,11),
TO_SIGNED(-77,11),
TO_SIGNED(-30,11),
TO_SIGNED(17,11),
TO_SIGNED(64,11),
TO_SIGNED(111,11),
TO_SIGNED(157,11),
TO_SIGNED(203,11),
TO_SIGNED(247,11),
TO_SIGNED(291,11),
TO_SIGNED(334,11),
TO_SIGNED(375,11),
TO_SIGNED(415,11),
TO_SIGNED(454,11),
TO_SIGNED(490,11),
TO_SIGNED(525,11),
TO_SIGNED(557,11),
TO_SIGNED(588,11),
TO_SIGNED(616,11),
TO_SIGNED(641,11),
TO_SIGNED(664,11),
TO_SIGNED(685,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(709,11),
TO_SIGNED(692,11),
TO_SIGNED(673,11),
TO_SIGNED(651,11),
TO_SIGNED(626,11),
TO_SIGNED(599,11),
TO_SIGNED(569,11),
TO_SIGNED(538,11),
TO_SIGNED(504,11),
TO_SIGNED(468,11),
TO_SIGNED(430,11),
TO_SIGNED(391,11),
TO_SIGNED(350,11),
TO_SIGNED(308,11),
TO_SIGNED(265,11),
TO_SIGNED(220,11),
TO_SIGNED(175,11),
TO_SIGNED(129,11),
TO_SIGNED(82,11),
TO_SIGNED(35,11),
TO_SIGNED(-12,11),
TO_SIGNED(-59,11),
TO_SIGNED(-105,11),
TO_SIGNED(-152,11),
TO_SIGNED(-197,11),
TO_SIGNED(-242,11),
TO_SIGNED(-286,11),
TO_SIGNED(-329,11),
TO_SIGNED(-371,11),
TO_SIGNED(-411,11),
TO_SIGNED(-449,11),
TO_SIGNED(-486,11),
TO_SIGNED(-521,11),
TO_SIGNED(-554,11),
TO_SIGNED(-584,11),
TO_SIGNED(-613,11),
TO_SIGNED(-639,11),
TO_SIGNED(-662,11),
TO_SIGNED(-683,11),
TO_SIGNED(-701,11),
TO_SIGNED(-716,11),
TO_SIGNED(-729,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-711,11),
TO_SIGNED(-694,11),
TO_SIGNED(-675,11),
TO_SIGNED(-653,11),
TO_SIGNED(-629,11),
TO_SIGNED(-602,11),
TO_SIGNED(-573,11),
TO_SIGNED(-541,11),
TO_SIGNED(-508,11),
TO_SIGNED(-472,11),
TO_SIGNED(-435,11),
TO_SIGNED(-396,11),
TO_SIGNED(-355,11),
TO_SIGNED(-313,11),
TO_SIGNED(-270,11),
TO_SIGNED(-225,11),
TO_SIGNED(-180,11),
TO_SIGNED(-134,11),
TO_SIGNED(-87,11),
TO_SIGNED(-41,11),
TO_SIGNED(6,11),
TO_SIGNED(53,11),
TO_SIGNED(100,11),
TO_SIGNED(147,11),
TO_SIGNED(192,11),
TO_SIGNED(237,11),
TO_SIGNED(281,11),
TO_SIGNED(324,11),
TO_SIGNED(366,11),
TO_SIGNED(406,11),
TO_SIGNED(445,11),
TO_SIGNED(482,11),
TO_SIGNED(517,11),
TO_SIGNED(550,11),
TO_SIGNED(581,11),
TO_SIGNED(610,11),
TO_SIGNED(636,11),
TO_SIGNED(659,11),
TO_SIGNED(681,11),
TO_SIGNED(699,11),
TO_SIGNED(715,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(712,11),
TO_SIGNED(696,11),
TO_SIGNED(677,11),
TO_SIGNED(656,11),
TO_SIGNED(632,11),
TO_SIGNED(605,11),
TO_SIGNED(576,11),
TO_SIGNED(545,11),
TO_SIGNED(512,11),
TO_SIGNED(476,11),
TO_SIGNED(439,11),
TO_SIGNED(400,11),
TO_SIGNED(360,11),
TO_SIGNED(318,11),
TO_SIGNED(275,11),
TO_SIGNED(230,11),
TO_SIGNED(185,11),
TO_SIGNED(139,11),
TO_SIGNED(93,11),
TO_SIGNED(46,11),
TO_SIGNED(-1,11),
TO_SIGNED(-48,11),
TO_SIGNED(-95,11),
TO_SIGNED(-141,11),
TO_SIGNED(-187,11),
TO_SIGNED(-232,11),
TO_SIGNED(-276,11),
TO_SIGNED(-320,11),
TO_SIGNED(-362,11),
TO_SIGNED(-402,11),
TO_SIGNED(-441,11),
TO_SIGNED(-478,11),
TO_SIGNED(-513,11),
TO_SIGNED(-547,11),
TO_SIGNED(-578,11),
TO_SIGNED(-606,11),
TO_SIGNED(-633,11),
TO_SIGNED(-657,11),
TO_SIGNED(-678,11),
TO_SIGNED(-697,11),
TO_SIGNED(-713,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-714,11),
TO_SIGNED(-698,11),
TO_SIGNED(-680,11),
TO_SIGNED(-658,11),
TO_SIGNED(-635,11),
TO_SIGNED(-608,11),
TO_SIGNED(-580,11),
TO_SIGNED(-549,11),
TO_SIGNED(-516,11),
TO_SIGNED(-480,11),
TO_SIGNED(-443,11),
TO_SIGNED(-405,11),
TO_SIGNED(-364,11),
TO_SIGNED(-323,11),
TO_SIGNED(-279,11),
TO_SIGNED(-235,11),
TO_SIGNED(-190,11),
TO_SIGNED(-144,11),
TO_SIGNED(-98,11),
TO_SIGNED(-51,11),
TO_SIGNED(-4,11),
TO_SIGNED(43,11),
TO_SIGNED(90,11),
TO_SIGNED(136,11),
TO_SIGNED(182,11),
TO_SIGNED(227,11),
TO_SIGNED(272,11),
TO_SIGNED(315,11),
TO_SIGNED(357,11),
TO_SIGNED(397,11),
TO_SIGNED(437,11),
TO_SIGNED(474,11),
TO_SIGNED(509,11),
TO_SIGNED(543,11),
TO_SIGNED(574,11),
TO_SIGNED(603,11),
TO_SIGNED(630,11),
TO_SIGNED(654,11),
TO_SIGNED(676,11),
TO_SIGNED(695,11),
TO_SIGNED(711,11),
TO_SIGNED(725,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(716,11),
TO_SIGNED(700,11),
TO_SIGNED(682,11),
TO_SIGNED(661,11),
TO_SIGNED(637,11),
TO_SIGNED(611,11),
TO_SIGNED(583,11),
TO_SIGNED(552,11),
TO_SIGNED(519,11),
TO_SIGNED(485,11),
TO_SIGNED(448,11),
TO_SIGNED(409,11),
TO_SIGNED(369,11),
TO_SIGNED(327,11),
TO_SIGNED(284,11),
TO_SIGNED(240,11),
TO_SIGNED(195,11),
TO_SIGNED(150,11),
TO_SIGNED(103,11),
TO_SIGNED(57,11),
TO_SIGNED(10,11),
TO_SIGNED(-37,11),
TO_SIGNED(-84,11),
TO_SIGNED(-131,11),
TO_SIGNED(-177,11),
TO_SIGNED(-222,11),
TO_SIGNED(-267,11),
TO_SIGNED(-310,11),
TO_SIGNED(-352,11),
TO_SIGNED(-393,11),
TO_SIGNED(-432,11),
TO_SIGNED(-470,11),
TO_SIGNED(-505,11),
TO_SIGNED(-539,11),
TO_SIGNED(-571,11),
TO_SIGNED(-600,11),
TO_SIGNED(-627,11),
TO_SIGNED(-652,11),
TO_SIGNED(-674,11),
TO_SIGNED(-693,11),
TO_SIGNED(-710,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-702,11),
TO_SIGNED(-684,11),
TO_SIGNED(-663,11),
TO_SIGNED(-640,11),
TO_SIGNED(-615,11),
TO_SIGNED(-586,11),
TO_SIGNED(-556,11),
TO_SIGNED(-523,11),
TO_SIGNED(-489,11),
TO_SIGNED(-452,11),
TO_SIGNED(-414,11),
TO_SIGNED(-374,11),
TO_SIGNED(-332,11),
TO_SIGNED(-289,11),
TO_SIGNED(-245,11),
TO_SIGNED(-201,11),
TO_SIGNED(-155,11),
TO_SIGNED(-109,11),
TO_SIGNED(-62,11),
TO_SIGNED(-15,11),
TO_SIGNED(32,11),
TO_SIGNED(79,11),
TO_SIGNED(125,11),
TO_SIGNED(172,11),
TO_SIGNED(217,11),
TO_SIGNED(262,11),
TO_SIGNED(305,11),
TO_SIGNED(347,11),
TO_SIGNED(388,11),
TO_SIGNED(428,11),
TO_SIGNED(466,11),
TO_SIGNED(501,11),
TO_SIGNED(535,11),
TO_SIGNED(567,11),
TO_SIGNED(597,11),
TO_SIGNED(624,11),
TO_SIGNED(649,11),
TO_SIGNED(671,11),
TO_SIGNED(691,11),
TO_SIGNED(708,11),
TO_SIGNED(722,11),
TO_SIGNED(733,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(704,11),
TO_SIGNED(686,11),
TO_SIGNED(666,11),
TO_SIGNED(643,11),
TO_SIGNED(618,11),
TO_SIGNED(590,11),
TO_SIGNED(559,11),
TO_SIGNED(527,11),
TO_SIGNED(493,11),
TO_SIGNED(456,11),
TO_SIGNED(418,11),
TO_SIGNED(378,11),
TO_SIGNED(337,11),
TO_SIGNED(294,11),
TO_SIGNED(250,11),
TO_SIGNED(206,11),
TO_SIGNED(160,11),
TO_SIGNED(114,11),
TO_SIGNED(67,11),
TO_SIGNED(20,11),
TO_SIGNED(-27,11),
TO_SIGNED(-74,11),
TO_SIGNED(-120,11),
TO_SIGNED(-166,11),
TO_SIGNED(-212,11),
TO_SIGNED(-257,11),
TO_SIGNED(-300,11),
TO_SIGNED(-343,11),
TO_SIGNED(-384,11),
TO_SIGNED(-423,11),
TO_SIGNED(-461,11),
TO_SIGNED(-497,11),
TO_SIGNED(-532,11),
TO_SIGNED(-564,11),
TO_SIGNED(-594,11),
TO_SIGNED(-621,11),
TO_SIGNED(-646,11),
TO_SIGNED(-669,11),
TO_SIGNED(-689,11),
TO_SIGNED(-706,11),
TO_SIGNED(-721,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-720,11),
TO_SIGNED(-706,11),
TO_SIGNED(-688,11),
TO_SIGNED(-668,11),
TO_SIGNED(-646,11),
TO_SIGNED(-621,11),
TO_SIGNED(-593,11),
TO_SIGNED(-563,11),
TO_SIGNED(-531,11),
TO_SIGNED(-497,11),
TO_SIGNED(-460,11),
TO_SIGNED(-422,11),
TO_SIGNED(-383,11),
TO_SIGNED(-342,11),
TO_SIGNED(-299,11),
TO_SIGNED(-256,11),
TO_SIGNED(-211,11),
TO_SIGNED(-165,11),
TO_SIGNED(-119,11),
TO_SIGNED(-73,11),
TO_SIGNED(-26,11),
TO_SIGNED(21,11),
TO_SIGNED(68,11),
TO_SIGNED(115,11),
TO_SIGNED(161,11),
TO_SIGNED(207,11),
TO_SIGNED(251,11),
TO_SIGNED(295,11),
TO_SIGNED(338,11),
TO_SIGNED(379,11),
TO_SIGNED(419,11),
TO_SIGNED(457,11),
TO_SIGNED(493,11),
TO_SIGNED(528,11),
TO_SIGNED(560,11),
TO_SIGNED(590,11),
TO_SIGNED(618,11),
TO_SIGNED(644,11),
TO_SIGNED(666,11),
TO_SIGNED(687,11),
TO_SIGNED(704,11),
TO_SIGNED(719,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(671,11),
TO_SIGNED(648,11),
TO_SIGNED(624,11),
TO_SIGNED(596,11),
TO_SIGNED(567,11),
TO_SIGNED(535,11),
TO_SIGNED(501,11),
TO_SIGNED(465,11),
TO_SIGNED(427,11),
TO_SIGNED(387,11),
TO_SIGNED(346,11),
TO_SIGNED(304,11),
TO_SIGNED(261,11),
TO_SIGNED(216,11),
TO_SIGNED(171,11),
TO_SIGNED(124,11),
TO_SIGNED(78,11),
TO_SIGNED(31,11),
TO_SIGNED(-16,11),
TO_SIGNED(-63,11),
TO_SIGNED(-110,11),
TO_SIGNED(-156,11),
TO_SIGNED(-202,11),
TO_SIGNED(-246,11),
TO_SIGNED(-290,11),
TO_SIGNED(-333,11),
TO_SIGNED(-375,11),
TO_SIGNED(-415,11),
TO_SIGNED(-453,11),
TO_SIGNED(-489,11),
TO_SIGNED(-524,11),
TO_SIGNED(-557,11),
TO_SIGNED(-587,11),
TO_SIGNED(-615,11),
TO_SIGNED(-641,11),
TO_SIGNED(-664,11),
TO_SIGNED(-685,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-730,11),
TO_SIGNED(-739,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-693,11),
TO_SIGNED(-673,11),
TO_SIGNED(-651,11),
TO_SIGNED(-627,11),
TO_SIGNED(-599,11),
TO_SIGNED(-570,11),
TO_SIGNED(-538,11),
TO_SIGNED(-505,11),
TO_SIGNED(-469,11),
TO_SIGNED(-431,11),
TO_SIGNED(-392,11),
TO_SIGNED(-351,11),
TO_SIGNED(-309,11),
TO_SIGNED(-266,11),
TO_SIGNED(-221,11),
TO_SIGNED(-176,11),
TO_SIGNED(-130,11),
TO_SIGNED(-83,11),
TO_SIGNED(-36,11),
TO_SIGNED(11,11),
TO_SIGNED(58,11),
TO_SIGNED(104,11),
TO_SIGNED(151,11),
TO_SIGNED(196,11),
TO_SIGNED(241,11),
TO_SIGNED(285,11),
TO_SIGNED(328,11),
TO_SIGNED(370,11),
TO_SIGNED(410,11),
TO_SIGNED(449,11),
TO_SIGNED(485,11),
TO_SIGNED(520,11),
TO_SIGNED(553,11),
TO_SIGNED(584,11),
TO_SIGNED(612,11),
TO_SIGNED(638,11),
TO_SIGNED(661,11),
TO_SIGNED(682,11),
TO_SIGNED(700,11),
TO_SIGNED(716,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(725,11),
TO_SIGNED(711,11),
TO_SIGNED(695,11),
TO_SIGNED(675,11),
TO_SIGNED(654,11),
TO_SIGNED(629,11),
TO_SIGNED(603,11),
TO_SIGNED(574,11),
TO_SIGNED(542,11),
TO_SIGNED(509,11),
TO_SIGNED(473,11),
TO_SIGNED(436,11),
TO_SIGNED(397,11),
TO_SIGNED(356,11),
TO_SIGNED(314,11),
TO_SIGNED(271,11),
TO_SIGNED(226,11),
TO_SIGNED(181,11),
TO_SIGNED(135,11),
TO_SIGNED(88,11),
TO_SIGNED(42,11),
TO_SIGNED(-5,11),
TO_SIGNED(-52,11),
TO_SIGNED(-99,11),
TO_SIGNED(-145,11),
TO_SIGNED(-191,11),
TO_SIGNED(-236,11),
TO_SIGNED(-280,11),
TO_SIGNED(-323,11),
TO_SIGNED(-365,11),
TO_SIGNED(-406,11),
TO_SIGNED(-444,11),
TO_SIGNED(-481,11),
TO_SIGNED(-516,11),
TO_SIGNED(-549,11),
TO_SIGNED(-580,11),
TO_SIGNED(-609,11),
TO_SIGNED(-635,11),
TO_SIGNED(-659,11),
TO_SIGNED(-680,11),
TO_SIGNED(-699,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-736,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-678,11),
TO_SIGNED(-656,11),
TO_SIGNED(-632,11),
TO_SIGNED(-606,11),
TO_SIGNED(-577,11),
TO_SIGNED(-546,11),
TO_SIGNED(-512,11),
TO_SIGNED(-477,11),
TO_SIGNED(-440,11),
TO_SIGNED(-401,11),
TO_SIGNED(-361,11),
TO_SIGNED(-319,11),
TO_SIGNED(-275,11),
TO_SIGNED(-231,11),
TO_SIGNED(-186,11),
TO_SIGNED(-140,11),
TO_SIGNED(-94,11),
TO_SIGNED(-47,11),
TO_SIGNED(0,11),
TO_SIGNED(47,11),
TO_SIGNED(94,11),
TO_SIGNED(140,11),
TO_SIGNED(186,11),
TO_SIGNED(231,11),
TO_SIGNED(275,11),
TO_SIGNED(319,11),
TO_SIGNED(361,11),
TO_SIGNED(401,11),
TO_SIGNED(440,11),
TO_SIGNED(477,11),
TO_SIGNED(512,11),
TO_SIGNED(546,11),
TO_SIGNED(577,11),
TO_SIGNED(606,11),
TO_SIGNED(632,11),
TO_SIGNED(656,11),
TO_SIGNED(678,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(736,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(699,11),
TO_SIGNED(680,11),
TO_SIGNED(659,11),
TO_SIGNED(635,11),
TO_SIGNED(609,11),
TO_SIGNED(580,11),
TO_SIGNED(549,11),
TO_SIGNED(516,11),
TO_SIGNED(481,11),
TO_SIGNED(444,11),
TO_SIGNED(406,11),
TO_SIGNED(365,11),
TO_SIGNED(323,11),
TO_SIGNED(280,11),
TO_SIGNED(236,11),
TO_SIGNED(191,11),
TO_SIGNED(145,11),
TO_SIGNED(99,11),
TO_SIGNED(52,11),
TO_SIGNED(5,11),
TO_SIGNED(-42,11),
TO_SIGNED(-88,11),
TO_SIGNED(-135,11),
TO_SIGNED(-181,11),
TO_SIGNED(-226,11),
TO_SIGNED(-271,11),
TO_SIGNED(-314,11),
TO_SIGNED(-356,11),
TO_SIGNED(-397,11),
TO_SIGNED(-436,11),
TO_SIGNED(-473,11),
TO_SIGNED(-509,11),
TO_SIGNED(-542,11),
TO_SIGNED(-574,11),
TO_SIGNED(-603,11),
TO_SIGNED(-629,11),
TO_SIGNED(-654,11),
TO_SIGNED(-675,11),
TO_SIGNED(-695,11),
TO_SIGNED(-711,11),
TO_SIGNED(-725,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-716,11),
TO_SIGNED(-700,11),
TO_SIGNED(-682,11),
TO_SIGNED(-661,11),
TO_SIGNED(-638,11),
TO_SIGNED(-612,11),
TO_SIGNED(-584,11),
TO_SIGNED(-553,11),
TO_SIGNED(-520,11),
TO_SIGNED(-485,11),
TO_SIGNED(-449,11),
TO_SIGNED(-410,11),
TO_SIGNED(-370,11),
TO_SIGNED(-328,11),
TO_SIGNED(-285,11),
TO_SIGNED(-241,11),
TO_SIGNED(-196,11),
TO_SIGNED(-151,11),
TO_SIGNED(-104,11),
TO_SIGNED(-58,11),
TO_SIGNED(-11,11),
TO_SIGNED(36,11),
TO_SIGNED(83,11),
TO_SIGNED(130,11),
TO_SIGNED(176,11),
TO_SIGNED(221,11),
TO_SIGNED(266,11),
TO_SIGNED(309,11),
TO_SIGNED(351,11),
TO_SIGNED(392,11),
TO_SIGNED(431,11),
TO_SIGNED(469,11),
TO_SIGNED(505,11),
TO_SIGNED(538,11),
TO_SIGNED(570,11),
TO_SIGNED(599,11),
TO_SIGNED(627,11),
TO_SIGNED(651,11),
TO_SIGNED(673,11),
TO_SIGNED(693,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(739,11),
TO_SIGNED(730,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(685,11),
TO_SIGNED(664,11),
TO_SIGNED(641,11),
TO_SIGNED(615,11),
TO_SIGNED(587,11),
TO_SIGNED(557,11),
TO_SIGNED(524,11),
TO_SIGNED(489,11),
TO_SIGNED(453,11),
TO_SIGNED(415,11),
TO_SIGNED(375,11),
TO_SIGNED(333,11),
TO_SIGNED(290,11),
TO_SIGNED(246,11),
TO_SIGNED(202,11),
TO_SIGNED(156,11),
TO_SIGNED(110,11),
TO_SIGNED(63,11),
TO_SIGNED(16,11),
TO_SIGNED(-31,11),
TO_SIGNED(-78,11),
TO_SIGNED(-124,11),
TO_SIGNED(-171,11),
TO_SIGNED(-216,11),
TO_SIGNED(-261,11),
TO_SIGNED(-304,11),
TO_SIGNED(-346,11),
TO_SIGNED(-387,11),
TO_SIGNED(-427,11),
TO_SIGNED(-465,11),
TO_SIGNED(-501,11),
TO_SIGNED(-535,11),
TO_SIGNED(-567,11),
TO_SIGNED(-596,11),
TO_SIGNED(-624,11),
TO_SIGNED(-648,11),
TO_SIGNED(-671,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-719,11),
TO_SIGNED(-704,11),
TO_SIGNED(-687,11),
TO_SIGNED(-666,11),
TO_SIGNED(-644,11),
TO_SIGNED(-618,11),
TO_SIGNED(-590,11),
TO_SIGNED(-560,11),
TO_SIGNED(-528,11),
TO_SIGNED(-493,11),
TO_SIGNED(-457,11),
TO_SIGNED(-419,11),
TO_SIGNED(-379,11),
TO_SIGNED(-338,11),
TO_SIGNED(-295,11),
TO_SIGNED(-251,11),
TO_SIGNED(-207,11),
TO_SIGNED(-161,11),
TO_SIGNED(-115,11),
TO_SIGNED(-68,11),
TO_SIGNED(-21,11),
TO_SIGNED(26,11),
TO_SIGNED(73,11),
TO_SIGNED(119,11),
TO_SIGNED(165,11),
TO_SIGNED(211,11),
TO_SIGNED(256,11),
TO_SIGNED(299,11),
TO_SIGNED(342,11),
TO_SIGNED(383,11),
TO_SIGNED(422,11),
TO_SIGNED(460,11),
TO_SIGNED(497,11),
TO_SIGNED(531,11),
TO_SIGNED(563,11),
TO_SIGNED(593,11),
TO_SIGNED(621,11),
TO_SIGNED(646,11),
TO_SIGNED(668,11),
TO_SIGNED(688,11),
TO_SIGNED(706,11),
TO_SIGNED(720,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(721,11),
TO_SIGNED(706,11),
TO_SIGNED(689,11),
TO_SIGNED(669,11),
TO_SIGNED(646,11),
TO_SIGNED(621,11),
TO_SIGNED(594,11),
TO_SIGNED(564,11),
TO_SIGNED(532,11),
TO_SIGNED(497,11),
TO_SIGNED(461,11),
TO_SIGNED(423,11),
TO_SIGNED(384,11),
TO_SIGNED(343,11),
TO_SIGNED(300,11),
TO_SIGNED(257,11),
TO_SIGNED(212,11),
TO_SIGNED(166,11),
TO_SIGNED(120,11),
TO_SIGNED(74,11),
TO_SIGNED(27,11),
TO_SIGNED(-20,11),
TO_SIGNED(-67,11),
TO_SIGNED(-114,11),
TO_SIGNED(-160,11),
TO_SIGNED(-206,11),
TO_SIGNED(-250,11),
TO_SIGNED(-294,11),
TO_SIGNED(-337,11),
TO_SIGNED(-378,11),
TO_SIGNED(-418,11),
TO_SIGNED(-456,11),
TO_SIGNED(-493,11),
TO_SIGNED(-527,11),
TO_SIGNED(-559,11),
TO_SIGNED(-590,11),
TO_SIGNED(-618,11),
TO_SIGNED(-643,11),
TO_SIGNED(-666,11),
TO_SIGNED(-686,11),
TO_SIGNED(-704,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-733,11),
TO_SIGNED(-722,11),
TO_SIGNED(-708,11),
TO_SIGNED(-691,11),
TO_SIGNED(-671,11),
TO_SIGNED(-649,11),
TO_SIGNED(-624,11),
TO_SIGNED(-597,11),
TO_SIGNED(-567,11),
TO_SIGNED(-535,11),
TO_SIGNED(-501,11),
TO_SIGNED(-466,11),
TO_SIGNED(-428,11),
TO_SIGNED(-388,11),
TO_SIGNED(-347,11),
TO_SIGNED(-305,11),
TO_SIGNED(-262,11),
TO_SIGNED(-217,11),
TO_SIGNED(-172,11),
TO_SIGNED(-125,11),
TO_SIGNED(-79,11),
TO_SIGNED(-32,11),
TO_SIGNED(15,11),
TO_SIGNED(62,11),
TO_SIGNED(109,11),
TO_SIGNED(155,11),
TO_SIGNED(201,11),
TO_SIGNED(245,11),
TO_SIGNED(289,11),
TO_SIGNED(332,11),
TO_SIGNED(374,11),
TO_SIGNED(414,11),
TO_SIGNED(452,11),
TO_SIGNED(489,11),
TO_SIGNED(523,11),
TO_SIGNED(556,11),
TO_SIGNED(586,11),
TO_SIGNED(615,11),
TO_SIGNED(640,11),
TO_SIGNED(663,11),
TO_SIGNED(684,11),
TO_SIGNED(702,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(710,11),
TO_SIGNED(693,11),
TO_SIGNED(674,11),
TO_SIGNED(652,11),
TO_SIGNED(627,11),
TO_SIGNED(600,11),
TO_SIGNED(571,11),
TO_SIGNED(539,11),
TO_SIGNED(505,11),
TO_SIGNED(470,11),
TO_SIGNED(432,11),
TO_SIGNED(393,11),
TO_SIGNED(352,11),
TO_SIGNED(310,11),
TO_SIGNED(267,11),
TO_SIGNED(222,11),
TO_SIGNED(177,11),
TO_SIGNED(131,11),
TO_SIGNED(84,11),
TO_SIGNED(37,11),
TO_SIGNED(-10,11),
TO_SIGNED(-57,11),
TO_SIGNED(-103,11),
TO_SIGNED(-150,11),
TO_SIGNED(-195,11),
TO_SIGNED(-240,11),
TO_SIGNED(-284,11),
TO_SIGNED(-327,11),
TO_SIGNED(-369,11),
TO_SIGNED(-409,11),
TO_SIGNED(-448,11),
TO_SIGNED(-485,11),
TO_SIGNED(-519,11),
TO_SIGNED(-552,11),
TO_SIGNED(-583,11),
TO_SIGNED(-611,11),
TO_SIGNED(-637,11),
TO_SIGNED(-661,11),
TO_SIGNED(-682,11),
TO_SIGNED(-700,11),
TO_SIGNED(-716,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-725,11),
TO_SIGNED(-711,11),
TO_SIGNED(-695,11),
TO_SIGNED(-676,11),
TO_SIGNED(-654,11),
TO_SIGNED(-630,11),
TO_SIGNED(-603,11),
TO_SIGNED(-574,11),
TO_SIGNED(-543,11),
TO_SIGNED(-509,11),
TO_SIGNED(-474,11),
TO_SIGNED(-437,11),
TO_SIGNED(-397,11),
TO_SIGNED(-357,11),
TO_SIGNED(-315,11),
TO_SIGNED(-272,11),
TO_SIGNED(-227,11),
TO_SIGNED(-182,11),
TO_SIGNED(-136,11),
TO_SIGNED(-90,11),
TO_SIGNED(-43,11),
TO_SIGNED(4,11),
TO_SIGNED(51,11),
TO_SIGNED(98,11),
TO_SIGNED(144,11),
TO_SIGNED(190,11),
TO_SIGNED(235,11),
TO_SIGNED(279,11),
TO_SIGNED(323,11),
TO_SIGNED(364,11),
TO_SIGNED(405,11),
TO_SIGNED(443,11),
TO_SIGNED(480,11),
TO_SIGNED(516,11),
TO_SIGNED(549,11),
TO_SIGNED(580,11),
TO_SIGNED(608,11),
TO_SIGNED(635,11),
TO_SIGNED(658,11),
TO_SIGNED(680,11),
TO_SIGNED(698,11),
TO_SIGNED(714,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(713,11),
TO_SIGNED(697,11),
TO_SIGNED(678,11),
TO_SIGNED(657,11),
TO_SIGNED(633,11),
TO_SIGNED(606,11),
TO_SIGNED(578,11),
TO_SIGNED(547,11),
TO_SIGNED(513,11),
TO_SIGNED(478,11),
TO_SIGNED(441,11),
TO_SIGNED(402,11),
TO_SIGNED(362,11),
TO_SIGNED(320,11),
TO_SIGNED(276,11),
TO_SIGNED(232,11),
TO_SIGNED(187,11),
TO_SIGNED(141,11),
TO_SIGNED(95,11),
TO_SIGNED(48,11),
TO_SIGNED(1,11),
TO_SIGNED(-46,11),
TO_SIGNED(-93,11),
TO_SIGNED(-139,11),
TO_SIGNED(-185,11),
TO_SIGNED(-230,11),
TO_SIGNED(-275,11),
TO_SIGNED(-318,11),
TO_SIGNED(-360,11),
TO_SIGNED(-400,11),
TO_SIGNED(-439,11),
TO_SIGNED(-476,11),
TO_SIGNED(-512,11),
TO_SIGNED(-545,11),
TO_SIGNED(-576,11),
TO_SIGNED(-605,11),
TO_SIGNED(-632,11),
TO_SIGNED(-656,11),
TO_SIGNED(-677,11),
TO_SIGNED(-696,11),
TO_SIGNED(-712,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-715,11),
TO_SIGNED(-699,11),
TO_SIGNED(-681,11),
TO_SIGNED(-659,11),
TO_SIGNED(-636,11),
TO_SIGNED(-610,11),
TO_SIGNED(-581,11),
TO_SIGNED(-550,11),
TO_SIGNED(-517,11),
TO_SIGNED(-482,11),
TO_SIGNED(-445,11),
TO_SIGNED(-406,11),
TO_SIGNED(-366,11),
TO_SIGNED(-324,11),
TO_SIGNED(-281,11),
TO_SIGNED(-237,11),
TO_SIGNED(-192,11),
TO_SIGNED(-147,11),
TO_SIGNED(-100,11),
TO_SIGNED(-53,11),
TO_SIGNED(-6,11),
TO_SIGNED(41,11),
TO_SIGNED(87,11),
TO_SIGNED(134,11),
TO_SIGNED(180,11),
TO_SIGNED(225,11),
TO_SIGNED(270,11),
TO_SIGNED(313,11),
TO_SIGNED(355,11),
TO_SIGNED(396,11),
TO_SIGNED(435,11),
TO_SIGNED(472,11),
TO_SIGNED(508,11),
TO_SIGNED(541,11),
TO_SIGNED(573,11),
TO_SIGNED(602,11),
TO_SIGNED(629,11),
TO_SIGNED(653,11),
TO_SIGNED(675,11),
TO_SIGNED(694,11),
TO_SIGNED(711,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(729,11),
TO_SIGNED(716,11),
TO_SIGNED(701,11),
TO_SIGNED(683,11),
TO_SIGNED(662,11),
TO_SIGNED(639,11),
TO_SIGNED(613,11),
TO_SIGNED(584,11),
TO_SIGNED(554,11),
TO_SIGNED(521,11),
TO_SIGNED(486,11),
TO_SIGNED(449,11),
TO_SIGNED(411,11),
TO_SIGNED(371,11),
TO_SIGNED(329,11),
TO_SIGNED(286,11),
TO_SIGNED(242,11),
TO_SIGNED(197,11),
TO_SIGNED(152,11),
TO_SIGNED(105,11),
TO_SIGNED(59,11),
TO_SIGNED(12,11),
TO_SIGNED(-35,11),
TO_SIGNED(-82,11),
TO_SIGNED(-129,11),
TO_SIGNED(-175,11),
TO_SIGNED(-220,11),
TO_SIGNED(-265,11),
TO_SIGNED(-308,11),
TO_SIGNED(-350,11),
TO_SIGNED(-391,11),
TO_SIGNED(-430,11),
TO_SIGNED(-468,11),
TO_SIGNED(-504,11),
TO_SIGNED(-538,11),
TO_SIGNED(-569,11),
TO_SIGNED(-599,11),
TO_SIGNED(-626,11),
TO_SIGNED(-651,11),
TO_SIGNED(-673,11),
TO_SIGNED(-692,11),
TO_SIGNED(-709,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-685,11),
TO_SIGNED(-664,11),
TO_SIGNED(-641,11),
TO_SIGNED(-616,11),
TO_SIGNED(-588,11),
TO_SIGNED(-557,11),
TO_SIGNED(-525,11),
TO_SIGNED(-490,11),
TO_SIGNED(-454,11),
TO_SIGNED(-415,11),
TO_SIGNED(-375,11),
TO_SIGNED(-334,11),
TO_SIGNED(-291,11),
TO_SIGNED(-247,11),
TO_SIGNED(-203,11),
TO_SIGNED(-157,11),
TO_SIGNED(-111,11),
TO_SIGNED(-64,11),
TO_SIGNED(-17,11),
TO_SIGNED(30,11),
TO_SIGNED(77,11),
TO_SIGNED(123,11),
TO_SIGNED(169,11),
TO_SIGNED(215,11),
TO_SIGNED(260,11),
TO_SIGNED(303,11),
TO_SIGNED(345,11),
TO_SIGNED(387,11),
TO_SIGNED(426,11),
TO_SIGNED(464,11),
TO_SIGNED(500,11),
TO_SIGNED(534,11),
TO_SIGNED(566,11),
TO_SIGNED(596,11),
TO_SIGNED(623,11),
TO_SIGNED(648,11),
TO_SIGNED(670,11),
TO_SIGNED(690,11),
TO_SIGNED(707,11),
TO_SIGNED(721,11),
TO_SIGNED(733,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(705,11),
TO_SIGNED(687,11),
TO_SIGNED(667,11),
TO_SIGNED(644,11),
TO_SIGNED(619,11),
TO_SIGNED(591,11),
TO_SIGNED(561,11),
TO_SIGNED(529,11),
TO_SIGNED(494,11),
TO_SIGNED(458,11),
TO_SIGNED(420,11),
TO_SIGNED(380,11),
TO_SIGNED(339,11),
TO_SIGNED(296,11),
TO_SIGNED(252,11),
TO_SIGNED(208,11),
TO_SIGNED(162,11),
TO_SIGNED(116,11),
TO_SIGNED(69,11),
TO_SIGNED(22,11),
TO_SIGNED(-25,11),
TO_SIGNED(-71,11),
TO_SIGNED(-118,11),
TO_SIGNED(-164,11),
TO_SIGNED(-210,11),
TO_SIGNED(-255,11),
TO_SIGNED(-298,11),
TO_SIGNED(-341,11),
TO_SIGNED(-382,11),
TO_SIGNED(-422,11),
TO_SIGNED(-460,11),
TO_SIGNED(-496,11),
TO_SIGNED(-530,11),
TO_SIGNED(-562,11),
TO_SIGNED(-592,11),
TO_SIGNED(-620,11),
TO_SIGNED(-645,11),
TO_SIGNED(-668,11),
TO_SIGNED(-688,11),
TO_SIGNED(-705,11),
TO_SIGNED(-720,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-721,11),
TO_SIGNED(-706,11),
TO_SIGNED(-689,11),
TO_SIGNED(-669,11),
TO_SIGNED(-647,11),
TO_SIGNED(-622,11),
TO_SIGNED(-594,11),
TO_SIGNED(-564,11),
TO_SIGNED(-532,11),
TO_SIGNED(-498,11),
TO_SIGNED(-462,11),
TO_SIGNED(-424,11),
TO_SIGNED(-385,11),
TO_SIGNED(-344,11),
TO_SIGNED(-301,11),
TO_SIGNED(-258,11),
TO_SIGNED(-213,11),
TO_SIGNED(-167,11),
TO_SIGNED(-121,11),
TO_SIGNED(-75,11),
TO_SIGNED(-28,11),
TO_SIGNED(19,11),
TO_SIGNED(66,11),
TO_SIGNED(113,11),
TO_SIGNED(159,11),
TO_SIGNED(205,11),
TO_SIGNED(249,11),
TO_SIGNED(293,11),
TO_SIGNED(336,11),
TO_SIGNED(377,11),
TO_SIGNED(417,11),
TO_SIGNED(455,11),
TO_SIGNED(492,11),
TO_SIGNED(526,11),
TO_SIGNED(559,11),
TO_SIGNED(589,11),
TO_SIGNED(617,11),
TO_SIGNED(642,11),
TO_SIGNED(665,11),
TO_SIGNED(686,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(708,11),
TO_SIGNED(691,11),
TO_SIGNED(672,11),
TO_SIGNED(650,11),
TO_SIGNED(625,11),
TO_SIGNED(598,11),
TO_SIGNED(568,11),
TO_SIGNED(536,11),
TO_SIGNED(502,11),
TO_SIGNED(466,11),
TO_SIGNED(429,11),
TO_SIGNED(389,11),
TO_SIGNED(348,11),
TO_SIGNED(306,11),
TO_SIGNED(263,11),
TO_SIGNED(218,11),
TO_SIGNED(173,11),
TO_SIGNED(127,11),
TO_SIGNED(80,11),
TO_SIGNED(33,11),
TO_SIGNED(-14,11),
TO_SIGNED(-61,11),
TO_SIGNED(-108,11),
TO_SIGNED(-154,11),
TO_SIGNED(-200,11),
TO_SIGNED(-244,11),
TO_SIGNED(-288,11),
TO_SIGNED(-331,11),
TO_SIGNED(-373,11),
TO_SIGNED(-413,11),
TO_SIGNED(-451,11),
TO_SIGNED(-488,11),
TO_SIGNED(-523,11),
TO_SIGNED(-555,11),
TO_SIGNED(-586,11),
TO_SIGNED(-614,11),
TO_SIGNED(-640,11),
TO_SIGNED(-663,11),
TO_SIGNED(-684,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-729,11),
TO_SIGNED(-739,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-710,11),
TO_SIGNED(-693,11),
TO_SIGNED(-674,11),
TO_SIGNED(-652,11),
TO_SIGNED(-628,11),
TO_SIGNED(-601,11),
TO_SIGNED(-571,11),
TO_SIGNED(-540,11),
TO_SIGNED(-506,11),
TO_SIGNED(-471,11),
TO_SIGNED(-433,11),
TO_SIGNED(-394,11),
TO_SIGNED(-353,11),
TO_SIGNED(-311,11),
TO_SIGNED(-268,11),
TO_SIGNED(-223,11),
TO_SIGNED(-178,11),
TO_SIGNED(-132,11),
TO_SIGNED(-85,11),
TO_SIGNED(-38,11),
TO_SIGNED(9,11),
TO_SIGNED(56,11),
TO_SIGNED(102,11),
TO_SIGNED(149,11),
TO_SIGNED(194,11),
TO_SIGNED(239,11),
TO_SIGNED(283,11),
TO_SIGNED(326,11),
TO_SIGNED(368,11),
TO_SIGNED(408,11),
TO_SIGNED(447,11),
TO_SIGNED(484,11),
TO_SIGNED(519,11),
TO_SIGNED(552,11),
TO_SIGNED(582,11),
TO_SIGNED(611,11),
TO_SIGNED(637,11),
TO_SIGNED(660,11),
TO_SIGNED(681,11),
TO_SIGNED(700,11),
TO_SIGNED(715,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(736,11),
TO_SIGNED(725,11),
TO_SIGNED(712,11),
TO_SIGNED(695,11),
TO_SIGNED(676,11),
TO_SIGNED(655,11),
TO_SIGNED(631,11),
TO_SIGNED(604,11),
TO_SIGNED(575,11),
TO_SIGNED(544,11),
TO_SIGNED(510,11),
TO_SIGNED(475,11),
TO_SIGNED(437,11),
TO_SIGNED(398,11),
TO_SIGNED(358,11),
TO_SIGNED(316,11),
TO_SIGNED(273,11),
TO_SIGNED(228,11),
TO_SIGNED(183,11),
TO_SIGNED(137,11),
TO_SIGNED(91,11),
TO_SIGNED(44,11),
TO_SIGNED(-3,11),
TO_SIGNED(-50,11),
TO_SIGNED(-97,11),
TO_SIGNED(-143,11),
TO_SIGNED(-189,11),
TO_SIGNED(-234,11),
TO_SIGNED(-278,11),
TO_SIGNED(-322,11),
TO_SIGNED(-363,11),
TO_SIGNED(-404,11),
TO_SIGNED(-443,11),
TO_SIGNED(-480,11),
TO_SIGNED(-515,11),
TO_SIGNED(-548,11),
TO_SIGNED(-579,11),
TO_SIGNED(-608,11),
TO_SIGNED(-634,11),
TO_SIGNED(-658,11),
TO_SIGNED(-679,11),
TO_SIGNED(-698,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-679,11),
TO_SIGNED(-657,11),
TO_SIGNED(-633,11),
TO_SIGNED(-607,11),
TO_SIGNED(-578,11),
TO_SIGNED(-547,11),
TO_SIGNED(-514,11),
TO_SIGNED(-479,11),
TO_SIGNED(-442,11),
TO_SIGNED(-403,11),
TO_SIGNED(-362,11),
TO_SIGNED(-321,11),
TO_SIGNED(-277,11),
TO_SIGNED(-233,11),
TO_SIGNED(-188,11),
TO_SIGNED(-142,11),
TO_SIGNED(-96,11),
TO_SIGNED(-49,11),
TO_SIGNED(-2,11),
TO_SIGNED(45,11),
TO_SIGNED(92,11),
TO_SIGNED(138,11),
TO_SIGNED(184,11),
TO_SIGNED(229,11),
TO_SIGNED(274,11),
TO_SIGNED(317,11),
TO_SIGNED(359,11),
TO_SIGNED(399,11),
TO_SIGNED(438,11),
TO_SIGNED(476,11),
TO_SIGNED(511,11),
TO_SIGNED(544,11),
TO_SIGNED(576,11),
TO_SIGNED(605,11),
TO_SIGNED(631,11),
TO_SIGNED(655,11),
TO_SIGNED(677,11),
TO_SIGNED(696,11),
TO_SIGNED(712,11),
TO_SIGNED(725,11),
TO_SIGNED(736,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(715,11),
TO_SIGNED(699,11),
TO_SIGNED(681,11),
TO_SIGNED(660,11),
TO_SIGNED(636,11),
TO_SIGNED(610,11),
TO_SIGNED(582,11),
TO_SIGNED(551,11),
TO_SIGNED(518,11),
TO_SIGNED(483,11),
TO_SIGNED(446,11),
TO_SIGNED(407,11),
TO_SIGNED(367,11),
TO_SIGNED(325,11),
TO_SIGNED(282,11),
TO_SIGNED(238,11),
TO_SIGNED(193,11),
TO_SIGNED(148,11),
TO_SIGNED(101,11),
TO_SIGNED(54,11),
TO_SIGNED(7,11),
TO_SIGNED(-40,11),
TO_SIGNED(-86,11),
TO_SIGNED(-133,11),
TO_SIGNED(-179,11),
TO_SIGNED(-224,11),
TO_SIGNED(-269,11),
TO_SIGNED(-312,11),
TO_SIGNED(-354,11),
TO_SIGNED(-395,11),
TO_SIGNED(-434,11),
TO_SIGNED(-471,11),
TO_SIGNED(-507,11),
TO_SIGNED(-541,11),
TO_SIGNED(-572,11),
TO_SIGNED(-601,11),
TO_SIGNED(-628,11),
TO_SIGNED(-653,11),
TO_SIGNED(-675,11),
TO_SIGNED(-694,11),
TO_SIGNED(-710,11),
TO_SIGNED(-724,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-701,11),
TO_SIGNED(-683,11),
TO_SIGNED(-662,11),
TO_SIGNED(-639,11),
TO_SIGNED(-613,11),
TO_SIGNED(-585,11),
TO_SIGNED(-554,11),
TO_SIGNED(-522,11),
TO_SIGNED(-487,11),
TO_SIGNED(-450,11),
TO_SIGNED(-412,11),
TO_SIGNED(-372,11),
TO_SIGNED(-330,11),
TO_SIGNED(-287,11),
TO_SIGNED(-243,11),
TO_SIGNED(-198,11),
TO_SIGNED(-153,11),
TO_SIGNED(-106,11),
TO_SIGNED(-60,11),
TO_SIGNED(-13,11),
TO_SIGNED(34,11),
TO_SIGNED(81,11),
TO_SIGNED(128,11),
TO_SIGNED(174,11),
TO_SIGNED(219,11),
TO_SIGNED(264,11),
TO_SIGNED(307,11),
TO_SIGNED(349,11),
TO_SIGNED(390,11),
TO_SIGNED(430,11),
TO_SIGNED(467,11),
TO_SIGNED(503,11),
TO_SIGNED(537,11),
TO_SIGNED(569,11),
TO_SIGNED(598,11),
TO_SIGNED(625,11),
TO_SIGNED(650,11),
TO_SIGNED(672,11),
TO_SIGNED(692,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(730,11),
TO_SIGNED(718,11),
TO_SIGNED(703,11),
TO_SIGNED(685,11),
TO_SIGNED(665,11),
TO_SIGNED(642,11),
TO_SIGNED(616,11),
TO_SIGNED(588,11),
TO_SIGNED(558,11),
TO_SIGNED(526,11),
TO_SIGNED(491,11),
TO_SIGNED(455,11),
TO_SIGNED(416,11),
TO_SIGNED(376,11),
TO_SIGNED(335,11),
TO_SIGNED(292,11),
TO_SIGNED(248,11),
TO_SIGNED(204,11),
TO_SIGNED(158,11),
TO_SIGNED(112,11),
TO_SIGNED(65,11),
TO_SIGNED(18,11),
TO_SIGNED(-29,11),
TO_SIGNED(-76,11),
TO_SIGNED(-122,11),
TO_SIGNED(-168,11),
TO_SIGNED(-214,11),
TO_SIGNED(-259,11),
TO_SIGNED(-302,11),
TO_SIGNED(-345,11),
TO_SIGNED(-386,11),
TO_SIGNED(-425,11),
TO_SIGNED(-463,11),
TO_SIGNED(-499,11),
TO_SIGNED(-533,11),
TO_SIGNED(-565,11),
TO_SIGNED(-595,11),
TO_SIGNED(-622,11),
TO_SIGNED(-647,11),
TO_SIGNED(-670,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-721,11),
TO_SIGNED(-733,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-720,11),
TO_SIGNED(-705,11),
TO_SIGNED(-688,11),
TO_SIGNED(-667,11),
TO_SIGNED(-645,11),
TO_SIGNED(-619,11),
TO_SIGNED(-592,11),
TO_SIGNED(-562,11),
TO_SIGNED(-529,11),
TO_SIGNED(-495,11),
TO_SIGNED(-459,11),
TO_SIGNED(-421,11),
TO_SIGNED(-381,11),
TO_SIGNED(-340,11),
TO_SIGNED(-297,11),
TO_SIGNED(-254,11),
TO_SIGNED(-209,11),
TO_SIGNED(-163,11),
TO_SIGNED(-117,11),
TO_SIGNED(-70,11),
TO_SIGNED(-24,11),
TO_SIGNED(24,11),
TO_SIGNED(70,11),
TO_SIGNED(117,11),
TO_SIGNED(163,11),
TO_SIGNED(209,11),
TO_SIGNED(254,11),
TO_SIGNED(297,11),
TO_SIGNED(340,11),
TO_SIGNED(381,11),
TO_SIGNED(421,11),
TO_SIGNED(459,11),
TO_SIGNED(495,11),
TO_SIGNED(529,11),
TO_SIGNED(562,11),
TO_SIGNED(592,11),
TO_SIGNED(619,11),
TO_SIGNED(645,11),
TO_SIGNED(667,11),
TO_SIGNED(688,11),
TO_SIGNED(705,11),
TO_SIGNED(720,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(733,11),
TO_SIGNED(721,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(670,11),
TO_SIGNED(647,11),
TO_SIGNED(622,11),
TO_SIGNED(595,11),
TO_SIGNED(565,11),
TO_SIGNED(533,11),
TO_SIGNED(499,11),
TO_SIGNED(463,11),
TO_SIGNED(425,11),
TO_SIGNED(386,11),
TO_SIGNED(345,11),
TO_SIGNED(302,11),
TO_SIGNED(259,11),
TO_SIGNED(214,11),
TO_SIGNED(168,11),
TO_SIGNED(122,11),
TO_SIGNED(76,11),
TO_SIGNED(29,11),
TO_SIGNED(-18,11),
TO_SIGNED(-65,11),
TO_SIGNED(-112,11),
TO_SIGNED(-158,11),
TO_SIGNED(-204,11),
TO_SIGNED(-248,11),
TO_SIGNED(-292,11),
TO_SIGNED(-335,11),
TO_SIGNED(-376,11),
TO_SIGNED(-416,11),
TO_SIGNED(-455,11),
TO_SIGNED(-491,11),
TO_SIGNED(-526,11),
TO_SIGNED(-558,11),
TO_SIGNED(-588,11),
TO_SIGNED(-616,11),
TO_SIGNED(-642,11),
TO_SIGNED(-665,11),
TO_SIGNED(-685,11),
TO_SIGNED(-703,11),
TO_SIGNED(-718,11),
TO_SIGNED(-730,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-692,11),
TO_SIGNED(-672,11),
TO_SIGNED(-650,11),
TO_SIGNED(-625,11),
TO_SIGNED(-598,11),
TO_SIGNED(-569,11),
TO_SIGNED(-537,11),
TO_SIGNED(-503,11),
TO_SIGNED(-467,11),
TO_SIGNED(-430,11),
TO_SIGNED(-390,11),
TO_SIGNED(-349,11),
TO_SIGNED(-307,11),
TO_SIGNED(-264,11),
TO_SIGNED(-219,11),
TO_SIGNED(-174,11),
TO_SIGNED(-128,11),
TO_SIGNED(-81,11),
TO_SIGNED(-34,11),
TO_SIGNED(13,11),
TO_SIGNED(60,11),
TO_SIGNED(106,11),
TO_SIGNED(153,11),
TO_SIGNED(198,11),
TO_SIGNED(243,11),
TO_SIGNED(287,11),
TO_SIGNED(330,11),
TO_SIGNED(372,11),
TO_SIGNED(412,11),
TO_SIGNED(450,11),
TO_SIGNED(487,11),
TO_SIGNED(522,11),
TO_SIGNED(554,11),
TO_SIGNED(585,11),
TO_SIGNED(613,11),
TO_SIGNED(639,11),
TO_SIGNED(662,11),
TO_SIGNED(683,11),
TO_SIGNED(701,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(724,11),
TO_SIGNED(710,11),
TO_SIGNED(694,11),
TO_SIGNED(675,11),
TO_SIGNED(653,11),
TO_SIGNED(628,11),
TO_SIGNED(601,11),
TO_SIGNED(572,11),
TO_SIGNED(541,11),
TO_SIGNED(507,11),
TO_SIGNED(471,11),
TO_SIGNED(434,11),
TO_SIGNED(395,11),
TO_SIGNED(354,11),
TO_SIGNED(312,11),
TO_SIGNED(269,11),
TO_SIGNED(224,11),
TO_SIGNED(179,11),
TO_SIGNED(133,11),
TO_SIGNED(86,11),
TO_SIGNED(40,11),
TO_SIGNED(-7,11),
TO_SIGNED(-54,11),
TO_SIGNED(-101,11),
TO_SIGNED(-148,11),
TO_SIGNED(-193,11),
TO_SIGNED(-238,11),
TO_SIGNED(-282,11),
TO_SIGNED(-325,11),
TO_SIGNED(-367,11),
TO_SIGNED(-407,11),
TO_SIGNED(-446,11),
TO_SIGNED(-483,11),
TO_SIGNED(-518,11),
TO_SIGNED(-551,11),
TO_SIGNED(-582,11),
TO_SIGNED(-610,11),
TO_SIGNED(-636,11),
TO_SIGNED(-660,11),
TO_SIGNED(-681,11),
TO_SIGNED(-699,11),
TO_SIGNED(-715,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-736,11),
TO_SIGNED(-725,11),
TO_SIGNED(-712,11),
TO_SIGNED(-696,11),
TO_SIGNED(-677,11),
TO_SIGNED(-655,11),
TO_SIGNED(-631,11),
TO_SIGNED(-605,11),
TO_SIGNED(-576,11),
TO_SIGNED(-544,11),
TO_SIGNED(-511,11),
TO_SIGNED(-476,11),
TO_SIGNED(-438,11),
TO_SIGNED(-399,11),
TO_SIGNED(-359,11),
TO_SIGNED(-317,11),
TO_SIGNED(-274,11),
TO_SIGNED(-229,11),
TO_SIGNED(-184,11),
TO_SIGNED(-138,11),
TO_SIGNED(-92,11),
TO_SIGNED(-45,11),
TO_SIGNED(2,11),
TO_SIGNED(49,11),
TO_SIGNED(96,11),
TO_SIGNED(142,11),
TO_SIGNED(188,11),
TO_SIGNED(233,11),
TO_SIGNED(277,11),
TO_SIGNED(321,11),
TO_SIGNED(362,11),
TO_SIGNED(403,11),
TO_SIGNED(442,11),
TO_SIGNED(479,11),
TO_SIGNED(514,11),
TO_SIGNED(547,11),
TO_SIGNED(578,11),
TO_SIGNED(607,11),
TO_SIGNED(633,11),
TO_SIGNED(657,11),
TO_SIGNED(679,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(698,11),
TO_SIGNED(679,11),
TO_SIGNED(658,11),
TO_SIGNED(634,11),
TO_SIGNED(608,11),
TO_SIGNED(579,11),
TO_SIGNED(548,11),
TO_SIGNED(515,11),
TO_SIGNED(480,11),
TO_SIGNED(443,11),
TO_SIGNED(404,11),
TO_SIGNED(363,11),
TO_SIGNED(322,11),
TO_SIGNED(278,11),
TO_SIGNED(234,11),
TO_SIGNED(189,11),
TO_SIGNED(143,11),
TO_SIGNED(97,11),
TO_SIGNED(50,11),
TO_SIGNED(3,11),
TO_SIGNED(-44,11),
TO_SIGNED(-91,11),
TO_SIGNED(-137,11),
TO_SIGNED(-183,11),
TO_SIGNED(-228,11),
TO_SIGNED(-273,11),
TO_SIGNED(-316,11),
TO_SIGNED(-358,11),
TO_SIGNED(-398,11),
TO_SIGNED(-437,11),
TO_SIGNED(-475,11),
TO_SIGNED(-510,11),
TO_SIGNED(-544,11),
TO_SIGNED(-575,11),
TO_SIGNED(-604,11),
TO_SIGNED(-631,11),
TO_SIGNED(-655,11),
TO_SIGNED(-676,11),
TO_SIGNED(-695,11),
TO_SIGNED(-712,11),
TO_SIGNED(-725,11),
TO_SIGNED(-736,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-715,11),
TO_SIGNED(-700,11),
TO_SIGNED(-681,11),
TO_SIGNED(-660,11),
TO_SIGNED(-637,11),
TO_SIGNED(-611,11),
TO_SIGNED(-582,11),
TO_SIGNED(-552,11),
TO_SIGNED(-519,11),
TO_SIGNED(-484,11),
TO_SIGNED(-447,11),
TO_SIGNED(-408,11),
TO_SIGNED(-368,11),
TO_SIGNED(-326,11),
TO_SIGNED(-283,11),
TO_SIGNED(-239,11),
TO_SIGNED(-194,11),
TO_SIGNED(-149,11),
TO_SIGNED(-102,11),
TO_SIGNED(-56,11),
TO_SIGNED(-9,11),
TO_SIGNED(38,11),
TO_SIGNED(85,11),
TO_SIGNED(132,11),
TO_SIGNED(178,11),
TO_SIGNED(223,11),
TO_SIGNED(268,11),
TO_SIGNED(311,11),
TO_SIGNED(353,11),
TO_SIGNED(394,11),
TO_SIGNED(433,11),
TO_SIGNED(471,11),
TO_SIGNED(506,11),
TO_SIGNED(540,11),
TO_SIGNED(571,11),
TO_SIGNED(601,11),
TO_SIGNED(628,11),
TO_SIGNED(652,11),
TO_SIGNED(674,11),
TO_SIGNED(693,11),
TO_SIGNED(710,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(739,11),
TO_SIGNED(729,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(684,11),
TO_SIGNED(663,11),
TO_SIGNED(640,11),
TO_SIGNED(614,11),
TO_SIGNED(586,11),
TO_SIGNED(555,11),
TO_SIGNED(523,11),
TO_SIGNED(488,11),
TO_SIGNED(451,11),
TO_SIGNED(413,11),
TO_SIGNED(373,11),
TO_SIGNED(331,11),
TO_SIGNED(288,11),
TO_SIGNED(244,11),
TO_SIGNED(200,11),
TO_SIGNED(154,11),
TO_SIGNED(108,11),
TO_SIGNED(61,11),
TO_SIGNED(14,11),
TO_SIGNED(-33,11),
TO_SIGNED(-80,11),
TO_SIGNED(-127,11),
TO_SIGNED(-173,11),
TO_SIGNED(-218,11),
TO_SIGNED(-263,11),
TO_SIGNED(-306,11),
TO_SIGNED(-348,11),
TO_SIGNED(-389,11),
TO_SIGNED(-429,11),
TO_SIGNED(-466,11),
TO_SIGNED(-502,11),
TO_SIGNED(-536,11),
TO_SIGNED(-568,11),
TO_SIGNED(-598,11),
TO_SIGNED(-625,11),
TO_SIGNED(-650,11),
TO_SIGNED(-672,11),
TO_SIGNED(-691,11),
TO_SIGNED(-708,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-686,11),
TO_SIGNED(-665,11),
TO_SIGNED(-642,11),
TO_SIGNED(-617,11),
TO_SIGNED(-589,11),
TO_SIGNED(-559,11),
TO_SIGNED(-526,11),
TO_SIGNED(-492,11),
TO_SIGNED(-455,11),
TO_SIGNED(-417,11),
TO_SIGNED(-377,11),
TO_SIGNED(-336,11),
TO_SIGNED(-293,11),
TO_SIGNED(-249,11),
TO_SIGNED(-205,11),
TO_SIGNED(-159,11),
TO_SIGNED(-113,11),
TO_SIGNED(-66,11),
TO_SIGNED(-19,11),
TO_SIGNED(28,11),
TO_SIGNED(75,11),
TO_SIGNED(121,11),
TO_SIGNED(167,11),
TO_SIGNED(213,11),
TO_SIGNED(258,11),
TO_SIGNED(301,11),
TO_SIGNED(344,11),
TO_SIGNED(385,11),
TO_SIGNED(424,11),
TO_SIGNED(462,11),
TO_SIGNED(498,11),
TO_SIGNED(532,11),
TO_SIGNED(564,11),
TO_SIGNED(594,11),
TO_SIGNED(622,11),
TO_SIGNED(647,11),
TO_SIGNED(669,11),
TO_SIGNED(689,11),
TO_SIGNED(706,11),
TO_SIGNED(721,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(720,11),
TO_SIGNED(705,11),
TO_SIGNED(688,11),
TO_SIGNED(668,11),
TO_SIGNED(645,11),
TO_SIGNED(620,11),
TO_SIGNED(592,11),
TO_SIGNED(562,11),
TO_SIGNED(530,11),
TO_SIGNED(496,11),
TO_SIGNED(460,11),
TO_SIGNED(422,11),
TO_SIGNED(382,11),
TO_SIGNED(341,11),
TO_SIGNED(298,11),
TO_SIGNED(255,11),
TO_SIGNED(210,11),
TO_SIGNED(164,11),
TO_SIGNED(118,11),
TO_SIGNED(71,11),
TO_SIGNED(25,11),
TO_SIGNED(-22,11),
TO_SIGNED(-69,11),
TO_SIGNED(-116,11),
TO_SIGNED(-162,11),
TO_SIGNED(-208,11),
TO_SIGNED(-252,11),
TO_SIGNED(-296,11),
TO_SIGNED(-339,11),
TO_SIGNED(-380,11),
TO_SIGNED(-420,11),
TO_SIGNED(-458,11),
TO_SIGNED(-494,11),
TO_SIGNED(-529,11),
TO_SIGNED(-561,11),
TO_SIGNED(-591,11),
TO_SIGNED(-619,11),
TO_SIGNED(-644,11),
TO_SIGNED(-667,11),
TO_SIGNED(-687,11),
TO_SIGNED(-705,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-733,11),
TO_SIGNED(-721,11),
TO_SIGNED(-707,11),
TO_SIGNED(-690,11),
TO_SIGNED(-670,11),
TO_SIGNED(-648,11),
TO_SIGNED(-623,11),
TO_SIGNED(-596,11),
TO_SIGNED(-566,11),
TO_SIGNED(-534,11),
TO_SIGNED(-500,11),
TO_SIGNED(-464,11),
TO_SIGNED(-426,11),
TO_SIGNED(-387,11),
TO_SIGNED(-345,11),
TO_SIGNED(-303,11),
TO_SIGNED(-260,11),
TO_SIGNED(-215,11),
TO_SIGNED(-169,11),
TO_SIGNED(-123,11),
TO_SIGNED(-77,11),
TO_SIGNED(-30,11),
TO_SIGNED(17,11),
TO_SIGNED(64,11),
TO_SIGNED(111,11),
TO_SIGNED(157,11),
TO_SIGNED(203,11),
TO_SIGNED(247,11),
TO_SIGNED(291,11),
TO_SIGNED(334,11),
TO_SIGNED(375,11),
TO_SIGNED(415,11),
TO_SIGNED(454,11),
TO_SIGNED(490,11),
TO_SIGNED(525,11),
TO_SIGNED(557,11),
TO_SIGNED(588,11),
TO_SIGNED(616,11),
TO_SIGNED(641,11),
TO_SIGNED(664,11),
TO_SIGNED(685,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(709,11),
TO_SIGNED(692,11),
TO_SIGNED(673,11),
TO_SIGNED(651,11),
TO_SIGNED(626,11),
TO_SIGNED(599,11),
TO_SIGNED(569,11),
TO_SIGNED(538,11),
TO_SIGNED(504,11),
TO_SIGNED(468,11),
TO_SIGNED(430,11),
TO_SIGNED(391,11),
TO_SIGNED(350,11),
TO_SIGNED(308,11),
TO_SIGNED(265,11),
TO_SIGNED(220,11),
TO_SIGNED(175,11),
TO_SIGNED(129,11),
TO_SIGNED(82,11),
TO_SIGNED(35,11),
TO_SIGNED(-12,11),
TO_SIGNED(-59,11),
TO_SIGNED(-105,11),
TO_SIGNED(-152,11),
TO_SIGNED(-197,11),
TO_SIGNED(-242,11),
TO_SIGNED(-286,11),
TO_SIGNED(-329,11),
TO_SIGNED(-371,11),
TO_SIGNED(-411,11),
TO_SIGNED(-449,11),
TO_SIGNED(-486,11),
TO_SIGNED(-521,11),
TO_SIGNED(-554,11),
TO_SIGNED(-584,11),
TO_SIGNED(-613,11),
TO_SIGNED(-639,11),
TO_SIGNED(-662,11),
TO_SIGNED(-683,11),
TO_SIGNED(-701,11),
TO_SIGNED(-716,11),
TO_SIGNED(-729,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-711,11),
TO_SIGNED(-694,11),
TO_SIGNED(-675,11),
TO_SIGNED(-653,11),
TO_SIGNED(-629,11),
TO_SIGNED(-602,11),
TO_SIGNED(-573,11),
TO_SIGNED(-541,11),
TO_SIGNED(-508,11),
TO_SIGNED(-472,11),
TO_SIGNED(-435,11),
TO_SIGNED(-396,11),
TO_SIGNED(-355,11),
TO_SIGNED(-313,11),
TO_SIGNED(-270,11),
TO_SIGNED(-225,11),
TO_SIGNED(-180,11),
TO_SIGNED(-134,11),
TO_SIGNED(-87,11),
TO_SIGNED(-41,11),
TO_SIGNED(6,11),
TO_SIGNED(53,11),
TO_SIGNED(100,11),
TO_SIGNED(147,11),
TO_SIGNED(192,11),
TO_SIGNED(237,11),
TO_SIGNED(281,11),
TO_SIGNED(324,11),
TO_SIGNED(366,11),
TO_SIGNED(406,11),
TO_SIGNED(445,11),
TO_SIGNED(482,11),
TO_SIGNED(517,11),
TO_SIGNED(550,11),
TO_SIGNED(581,11),
TO_SIGNED(610,11),
TO_SIGNED(636,11),
TO_SIGNED(659,11),
TO_SIGNED(681,11),
TO_SIGNED(699,11),
TO_SIGNED(715,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(712,11),
TO_SIGNED(696,11),
TO_SIGNED(677,11),
TO_SIGNED(656,11),
TO_SIGNED(632,11),
TO_SIGNED(605,11),
TO_SIGNED(576,11),
TO_SIGNED(545,11),
TO_SIGNED(512,11),
TO_SIGNED(476,11),
TO_SIGNED(439,11),
TO_SIGNED(400,11),
TO_SIGNED(360,11),
TO_SIGNED(318,11),
TO_SIGNED(275,11),
TO_SIGNED(230,11),
TO_SIGNED(185,11),
TO_SIGNED(139,11),
TO_SIGNED(93,11),
TO_SIGNED(46,11),
TO_SIGNED(-1,11),
TO_SIGNED(-48,11),
TO_SIGNED(-95,11),
TO_SIGNED(-141,11),
TO_SIGNED(-187,11),
TO_SIGNED(-232,11),
TO_SIGNED(-276,11),
TO_SIGNED(-320,11),
TO_SIGNED(-362,11),
TO_SIGNED(-402,11),
TO_SIGNED(-441,11),
TO_SIGNED(-478,11),
TO_SIGNED(-513,11),
TO_SIGNED(-547,11),
TO_SIGNED(-578,11),
TO_SIGNED(-606,11),
TO_SIGNED(-633,11),
TO_SIGNED(-657,11),
TO_SIGNED(-678,11),
TO_SIGNED(-697,11),
TO_SIGNED(-713,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-714,11),
TO_SIGNED(-698,11),
TO_SIGNED(-680,11),
TO_SIGNED(-658,11),
TO_SIGNED(-635,11),
TO_SIGNED(-608,11),
TO_SIGNED(-580,11),
TO_SIGNED(-549,11),
TO_SIGNED(-516,11),
TO_SIGNED(-480,11),
TO_SIGNED(-443,11),
TO_SIGNED(-405,11),
TO_SIGNED(-364,11),
TO_SIGNED(-323,11),
TO_SIGNED(-279,11),
TO_SIGNED(-235,11),
TO_SIGNED(-190,11),
TO_SIGNED(-144,11),
TO_SIGNED(-98,11),
TO_SIGNED(-51,11),
TO_SIGNED(-4,11),
TO_SIGNED(43,11),
TO_SIGNED(90,11),
TO_SIGNED(136,11),
TO_SIGNED(182,11),
TO_SIGNED(227,11),
TO_SIGNED(272,11),
TO_SIGNED(315,11),
TO_SIGNED(357,11),
TO_SIGNED(397,11),
TO_SIGNED(437,11),
TO_SIGNED(474,11),
TO_SIGNED(509,11),
TO_SIGNED(543,11),
TO_SIGNED(574,11),
TO_SIGNED(603,11),
TO_SIGNED(630,11),
TO_SIGNED(654,11),
TO_SIGNED(676,11),
TO_SIGNED(695,11),
TO_SIGNED(711,11),
TO_SIGNED(725,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(716,11),
TO_SIGNED(700,11),
TO_SIGNED(682,11),
TO_SIGNED(661,11),
TO_SIGNED(637,11),
TO_SIGNED(611,11),
TO_SIGNED(583,11),
TO_SIGNED(552,11),
TO_SIGNED(519,11),
TO_SIGNED(485,11),
TO_SIGNED(448,11),
TO_SIGNED(409,11),
TO_SIGNED(369,11),
TO_SIGNED(327,11),
TO_SIGNED(284,11),
TO_SIGNED(240,11),
TO_SIGNED(195,11),
TO_SIGNED(150,11),
TO_SIGNED(103,11),
TO_SIGNED(57,11),
TO_SIGNED(10,11),
TO_SIGNED(-37,11),
TO_SIGNED(-84,11),
TO_SIGNED(-131,11),
TO_SIGNED(-177,11),
TO_SIGNED(-222,11),
TO_SIGNED(-267,11),
TO_SIGNED(-310,11),
TO_SIGNED(-352,11),
TO_SIGNED(-393,11),
TO_SIGNED(-432,11),
TO_SIGNED(-470,11),
TO_SIGNED(-505,11),
TO_SIGNED(-539,11),
TO_SIGNED(-571,11),
TO_SIGNED(-600,11),
TO_SIGNED(-627,11),
TO_SIGNED(-652,11),
TO_SIGNED(-674,11),
TO_SIGNED(-693,11),
TO_SIGNED(-710,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-702,11),
TO_SIGNED(-684,11),
TO_SIGNED(-663,11),
TO_SIGNED(-640,11),
TO_SIGNED(-615,11),
TO_SIGNED(-586,11),
TO_SIGNED(-556,11),
TO_SIGNED(-523,11),
TO_SIGNED(-489,11),
TO_SIGNED(-452,11),
TO_SIGNED(-414,11),
TO_SIGNED(-374,11),
TO_SIGNED(-332,11),
TO_SIGNED(-289,11),
TO_SIGNED(-245,11),
TO_SIGNED(-201,11),
TO_SIGNED(-155,11),
TO_SIGNED(-109,11),
TO_SIGNED(-62,11),
TO_SIGNED(-15,11),
TO_SIGNED(32,11),
TO_SIGNED(79,11),
TO_SIGNED(125,11),
TO_SIGNED(172,11),
TO_SIGNED(217,11),
TO_SIGNED(262,11),
TO_SIGNED(305,11),
TO_SIGNED(347,11),
TO_SIGNED(388,11),
TO_SIGNED(428,11),
TO_SIGNED(466,11),
TO_SIGNED(501,11),
TO_SIGNED(535,11),
TO_SIGNED(567,11),
TO_SIGNED(597,11),
TO_SIGNED(624,11),
TO_SIGNED(649,11),
TO_SIGNED(671,11),
TO_SIGNED(691,11),
TO_SIGNED(708,11),
TO_SIGNED(722,11),
TO_SIGNED(733,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(704,11),
TO_SIGNED(686,11),
TO_SIGNED(666,11),
TO_SIGNED(643,11),
TO_SIGNED(618,11),
TO_SIGNED(590,11),
TO_SIGNED(559,11),
TO_SIGNED(527,11),
TO_SIGNED(493,11),
TO_SIGNED(456,11),
TO_SIGNED(418,11),
TO_SIGNED(378,11),
TO_SIGNED(337,11),
TO_SIGNED(294,11),
TO_SIGNED(250,11),
TO_SIGNED(206,11),
TO_SIGNED(160,11),
TO_SIGNED(114,11),
TO_SIGNED(67,11),
TO_SIGNED(20,11),
TO_SIGNED(-27,11),
TO_SIGNED(-74,11),
TO_SIGNED(-120,11),
TO_SIGNED(-166,11),
TO_SIGNED(-212,11),
TO_SIGNED(-257,11),
TO_SIGNED(-300,11),
TO_SIGNED(-343,11),
TO_SIGNED(-384,11),
TO_SIGNED(-423,11),
TO_SIGNED(-461,11),
TO_SIGNED(-497,11),
TO_SIGNED(-532,11),
TO_SIGNED(-564,11),
TO_SIGNED(-594,11),
TO_SIGNED(-621,11),
TO_SIGNED(-646,11),
TO_SIGNED(-669,11),
TO_SIGNED(-689,11),
TO_SIGNED(-706,11),
TO_SIGNED(-721,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-720,11),
TO_SIGNED(-706,11),
TO_SIGNED(-688,11),
TO_SIGNED(-668,11),
TO_SIGNED(-646,11),
TO_SIGNED(-621,11),
TO_SIGNED(-593,11),
TO_SIGNED(-563,11),
TO_SIGNED(-531,11),
TO_SIGNED(-497,11),
TO_SIGNED(-460,11),
TO_SIGNED(-422,11),
TO_SIGNED(-383,11),
TO_SIGNED(-342,11),
TO_SIGNED(-299,11),
TO_SIGNED(-256,11),
TO_SIGNED(-211,11),
TO_SIGNED(-165,11),
TO_SIGNED(-119,11),
TO_SIGNED(-73,11),
TO_SIGNED(-26,11),
TO_SIGNED(21,11),
TO_SIGNED(68,11),
TO_SIGNED(115,11),
TO_SIGNED(161,11),
TO_SIGNED(207,11),
TO_SIGNED(251,11),
TO_SIGNED(295,11),
TO_SIGNED(338,11),
TO_SIGNED(379,11),
TO_SIGNED(419,11),
TO_SIGNED(457,11),
TO_SIGNED(493,11),
TO_SIGNED(528,11),
TO_SIGNED(560,11),
TO_SIGNED(590,11),
TO_SIGNED(618,11),
TO_SIGNED(644,11),
TO_SIGNED(666,11),
TO_SIGNED(687,11),
TO_SIGNED(704,11),
TO_SIGNED(719,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(671,11),
TO_SIGNED(648,11),
TO_SIGNED(624,11),
TO_SIGNED(596,11),
TO_SIGNED(567,11),
TO_SIGNED(535,11),
TO_SIGNED(501,11),
TO_SIGNED(465,11),
TO_SIGNED(427,11),
TO_SIGNED(387,11),
TO_SIGNED(346,11),
TO_SIGNED(304,11),
TO_SIGNED(261,11),
TO_SIGNED(216,11),
TO_SIGNED(171,11),
TO_SIGNED(124,11),
TO_SIGNED(78,11),
TO_SIGNED(31,11),
TO_SIGNED(-16,11),
TO_SIGNED(-63,11),
TO_SIGNED(-110,11),
TO_SIGNED(-156,11),
TO_SIGNED(-202,11),
TO_SIGNED(-246,11),
TO_SIGNED(-290,11),
TO_SIGNED(-333,11),
TO_SIGNED(-375,11),
TO_SIGNED(-415,11),
TO_SIGNED(-453,11),
TO_SIGNED(-489,11),
TO_SIGNED(-524,11),
TO_SIGNED(-557,11),
TO_SIGNED(-587,11),
TO_SIGNED(-615,11),
TO_SIGNED(-641,11),
TO_SIGNED(-664,11),
TO_SIGNED(-685,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-730,11),
TO_SIGNED(-739,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-693,11),
TO_SIGNED(-673,11),
TO_SIGNED(-651,11),
TO_SIGNED(-627,11),
TO_SIGNED(-599,11),
TO_SIGNED(-570,11),
TO_SIGNED(-538,11),
TO_SIGNED(-505,11),
TO_SIGNED(-469,11),
TO_SIGNED(-431,11),
TO_SIGNED(-392,11),
TO_SIGNED(-351,11),
TO_SIGNED(-309,11),
TO_SIGNED(-266,11),
TO_SIGNED(-221,11),
TO_SIGNED(-176,11),
TO_SIGNED(-130,11),
TO_SIGNED(-83,11),
TO_SIGNED(-36,11),
TO_SIGNED(11,11),
TO_SIGNED(58,11),
TO_SIGNED(104,11),
TO_SIGNED(151,11),
TO_SIGNED(196,11),
TO_SIGNED(241,11),
TO_SIGNED(285,11),
TO_SIGNED(328,11),
TO_SIGNED(370,11),
TO_SIGNED(410,11),
TO_SIGNED(449,11),
TO_SIGNED(485,11),
TO_SIGNED(520,11),
TO_SIGNED(553,11),
TO_SIGNED(584,11),
TO_SIGNED(612,11),
TO_SIGNED(638,11),
TO_SIGNED(661,11),
TO_SIGNED(682,11),
TO_SIGNED(700,11),
TO_SIGNED(716,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(725,11),
TO_SIGNED(711,11),
TO_SIGNED(695,11),
TO_SIGNED(675,11),
TO_SIGNED(654,11),
TO_SIGNED(629,11),
TO_SIGNED(603,11),
TO_SIGNED(574,11),
TO_SIGNED(542,11),
TO_SIGNED(509,11),
TO_SIGNED(473,11),
TO_SIGNED(436,11),
TO_SIGNED(397,11),
TO_SIGNED(356,11),
TO_SIGNED(314,11),
TO_SIGNED(271,11),
TO_SIGNED(226,11),
TO_SIGNED(181,11),
TO_SIGNED(135,11),
TO_SIGNED(88,11),
TO_SIGNED(42,11),
TO_SIGNED(-5,11),
TO_SIGNED(-52,11),
TO_SIGNED(-99,11),
TO_SIGNED(-145,11),
TO_SIGNED(-191,11),
TO_SIGNED(-236,11),
TO_SIGNED(-280,11),
TO_SIGNED(-323,11),
TO_SIGNED(-365,11),
TO_SIGNED(-406,11),
TO_SIGNED(-444,11),
TO_SIGNED(-481,11),
TO_SIGNED(-516,11),
TO_SIGNED(-549,11),
TO_SIGNED(-580,11),
TO_SIGNED(-609,11),
TO_SIGNED(-635,11),
TO_SIGNED(-659,11),
TO_SIGNED(-680,11),
TO_SIGNED(-699,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-736,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-678,11),
TO_SIGNED(-656,11),
TO_SIGNED(-632,11),
TO_SIGNED(-606,11),
TO_SIGNED(-577,11),
TO_SIGNED(-546,11),
TO_SIGNED(-512,11),
TO_SIGNED(-477,11),
TO_SIGNED(-440,11),
TO_SIGNED(-401,11),
TO_SIGNED(-361,11),
TO_SIGNED(-319,11),
TO_SIGNED(-275,11),
TO_SIGNED(-231,11),
TO_SIGNED(-186,11),
TO_SIGNED(-140,11),
TO_SIGNED(-94,11),
TO_SIGNED(-47,11),
TO_SIGNED(0,11),
TO_SIGNED(47,11),
TO_SIGNED(94,11),
TO_SIGNED(140,11),
TO_SIGNED(186,11),
TO_SIGNED(231,11),
TO_SIGNED(275,11),
TO_SIGNED(319,11),
TO_SIGNED(361,11),
TO_SIGNED(401,11),
TO_SIGNED(440,11),
TO_SIGNED(477,11),
TO_SIGNED(512,11),
TO_SIGNED(546,11),
TO_SIGNED(577,11),
TO_SIGNED(606,11),
TO_SIGNED(632,11),
TO_SIGNED(656,11),
TO_SIGNED(678,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(736,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(699,11),
TO_SIGNED(680,11),
TO_SIGNED(659,11),
TO_SIGNED(635,11),
TO_SIGNED(609,11),
TO_SIGNED(580,11),
TO_SIGNED(549,11),
TO_SIGNED(516,11),
TO_SIGNED(481,11),
TO_SIGNED(444,11),
TO_SIGNED(406,11),
TO_SIGNED(365,11),
TO_SIGNED(323,11),
TO_SIGNED(280,11),
TO_SIGNED(236,11),
TO_SIGNED(191,11),
TO_SIGNED(145,11),
TO_SIGNED(99,11),
TO_SIGNED(52,11),
TO_SIGNED(5,11),
TO_SIGNED(-42,11),
TO_SIGNED(-88,11),
TO_SIGNED(-135,11),
TO_SIGNED(-181,11),
TO_SIGNED(-226,11),
TO_SIGNED(-271,11),
TO_SIGNED(-314,11),
TO_SIGNED(-356,11),
TO_SIGNED(-397,11),
TO_SIGNED(-436,11),
TO_SIGNED(-473,11),
TO_SIGNED(-509,11),
TO_SIGNED(-542,11),
TO_SIGNED(-574,11),
TO_SIGNED(-603,11),
TO_SIGNED(-629,11),
TO_SIGNED(-654,11),
TO_SIGNED(-675,11),
TO_SIGNED(-695,11),
TO_SIGNED(-711,11),
TO_SIGNED(-725,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-716,11),
TO_SIGNED(-700,11),
TO_SIGNED(-682,11),
TO_SIGNED(-661,11),
TO_SIGNED(-638,11),
TO_SIGNED(-612,11),
TO_SIGNED(-584,11),
TO_SIGNED(-553,11),
TO_SIGNED(-520,11),
TO_SIGNED(-485,11),
TO_SIGNED(-449,11),
TO_SIGNED(-410,11),
TO_SIGNED(-370,11),
TO_SIGNED(-328,11),
TO_SIGNED(-285,11),
TO_SIGNED(-241,11),
TO_SIGNED(-196,11),
TO_SIGNED(-151,11),
TO_SIGNED(-104,11),
TO_SIGNED(-58,11),
TO_SIGNED(-11,11),
TO_SIGNED(36,11),
TO_SIGNED(83,11),
TO_SIGNED(130,11),
TO_SIGNED(176,11),
TO_SIGNED(221,11),
TO_SIGNED(266,11),
TO_SIGNED(309,11),
TO_SIGNED(351,11),
TO_SIGNED(392,11),
TO_SIGNED(431,11),
TO_SIGNED(469,11),
TO_SIGNED(505,11),
TO_SIGNED(538,11),
TO_SIGNED(570,11),
TO_SIGNED(599,11),
TO_SIGNED(627,11),
TO_SIGNED(651,11),
TO_SIGNED(673,11),
TO_SIGNED(693,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(739,11),
TO_SIGNED(730,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(685,11),
TO_SIGNED(664,11),
TO_SIGNED(641,11),
TO_SIGNED(615,11),
TO_SIGNED(587,11),
TO_SIGNED(557,11),
TO_SIGNED(524,11),
TO_SIGNED(489,11),
TO_SIGNED(453,11),
TO_SIGNED(415,11),
TO_SIGNED(375,11),
TO_SIGNED(333,11),
TO_SIGNED(290,11),
TO_SIGNED(246,11),
TO_SIGNED(202,11),
TO_SIGNED(156,11),
TO_SIGNED(110,11),
TO_SIGNED(63,11),
TO_SIGNED(16,11),
TO_SIGNED(-31,11),
TO_SIGNED(-78,11),
TO_SIGNED(-124,11),
TO_SIGNED(-171,11),
TO_SIGNED(-216,11),
TO_SIGNED(-261,11),
TO_SIGNED(-304,11),
TO_SIGNED(-346,11),
TO_SIGNED(-387,11),
TO_SIGNED(-427,11),
TO_SIGNED(-465,11),
TO_SIGNED(-501,11),
TO_SIGNED(-535,11),
TO_SIGNED(-567,11),
TO_SIGNED(-596,11),
TO_SIGNED(-624,11),
TO_SIGNED(-648,11),
TO_SIGNED(-671,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-719,11),
TO_SIGNED(-704,11),
TO_SIGNED(-687,11),
TO_SIGNED(-666,11),
TO_SIGNED(-644,11),
TO_SIGNED(-618,11),
TO_SIGNED(-590,11),
TO_SIGNED(-560,11),
TO_SIGNED(-528,11),
TO_SIGNED(-493,11),
TO_SIGNED(-457,11),
TO_SIGNED(-419,11),
TO_SIGNED(-379,11),
TO_SIGNED(-338,11),
TO_SIGNED(-295,11),
TO_SIGNED(-251,11),
TO_SIGNED(-207,11),
TO_SIGNED(-161,11),
TO_SIGNED(-115,11),
TO_SIGNED(-68,11),
TO_SIGNED(-21,11),
TO_SIGNED(26,11),
TO_SIGNED(73,11),
TO_SIGNED(119,11),
TO_SIGNED(165,11),
TO_SIGNED(211,11),
TO_SIGNED(256,11),
TO_SIGNED(299,11),
TO_SIGNED(342,11),
TO_SIGNED(383,11),
TO_SIGNED(422,11),
TO_SIGNED(460,11),
TO_SIGNED(497,11),
TO_SIGNED(531,11),
TO_SIGNED(563,11),
TO_SIGNED(593,11),
TO_SIGNED(621,11),
TO_SIGNED(646,11),
TO_SIGNED(668,11),
TO_SIGNED(688,11),
TO_SIGNED(706,11),
TO_SIGNED(720,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(721,11),
TO_SIGNED(706,11),
TO_SIGNED(689,11),
TO_SIGNED(669,11),
TO_SIGNED(646,11),
TO_SIGNED(621,11),
TO_SIGNED(594,11),
TO_SIGNED(564,11),
TO_SIGNED(532,11),
TO_SIGNED(497,11),
TO_SIGNED(461,11),
TO_SIGNED(423,11),
TO_SIGNED(384,11),
TO_SIGNED(343,11),
TO_SIGNED(300,11),
TO_SIGNED(257,11),
TO_SIGNED(212,11),
TO_SIGNED(166,11),
TO_SIGNED(120,11),
TO_SIGNED(74,11),
TO_SIGNED(27,11),
TO_SIGNED(-20,11),
TO_SIGNED(-67,11),
TO_SIGNED(-114,11),
TO_SIGNED(-160,11),
TO_SIGNED(-206,11),
TO_SIGNED(-250,11),
TO_SIGNED(-294,11),
TO_SIGNED(-337,11),
TO_SIGNED(-378,11),
TO_SIGNED(-418,11),
TO_SIGNED(-456,11),
TO_SIGNED(-493,11),
TO_SIGNED(-527,11),
TO_SIGNED(-559,11),
TO_SIGNED(-590,11),
TO_SIGNED(-618,11),
TO_SIGNED(-643,11),
TO_SIGNED(-666,11),
TO_SIGNED(-686,11),
TO_SIGNED(-704,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-733,11),
TO_SIGNED(-722,11),
TO_SIGNED(-708,11),
TO_SIGNED(-691,11),
TO_SIGNED(-671,11),
TO_SIGNED(-649,11),
TO_SIGNED(-624,11),
TO_SIGNED(-597,11),
TO_SIGNED(-567,11),
TO_SIGNED(-535,11),
TO_SIGNED(-501,11),
TO_SIGNED(-466,11),
TO_SIGNED(-428,11),
TO_SIGNED(-388,11),
TO_SIGNED(-347,11),
TO_SIGNED(-305,11),
TO_SIGNED(-262,11),
TO_SIGNED(-217,11),
TO_SIGNED(-172,11),
TO_SIGNED(-125,11),
TO_SIGNED(-79,11),
TO_SIGNED(-32,11),
TO_SIGNED(15,11),
TO_SIGNED(62,11),
TO_SIGNED(109,11),
TO_SIGNED(155,11),
TO_SIGNED(201,11),
TO_SIGNED(245,11),
TO_SIGNED(289,11),
TO_SIGNED(332,11),
TO_SIGNED(374,11),
TO_SIGNED(414,11),
TO_SIGNED(452,11),
TO_SIGNED(489,11),
TO_SIGNED(523,11),
TO_SIGNED(556,11),
TO_SIGNED(586,11),
TO_SIGNED(615,11),
TO_SIGNED(640,11),
TO_SIGNED(663,11),
TO_SIGNED(684,11),
TO_SIGNED(702,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(710,11),
TO_SIGNED(693,11),
TO_SIGNED(674,11),
TO_SIGNED(652,11),
TO_SIGNED(627,11),
TO_SIGNED(600,11),
TO_SIGNED(571,11),
TO_SIGNED(539,11),
TO_SIGNED(505,11),
TO_SIGNED(470,11),
TO_SIGNED(432,11),
TO_SIGNED(393,11),
TO_SIGNED(352,11),
TO_SIGNED(310,11),
TO_SIGNED(267,11),
TO_SIGNED(222,11),
TO_SIGNED(177,11),
TO_SIGNED(131,11),
TO_SIGNED(84,11),
TO_SIGNED(37,11),
TO_SIGNED(-10,11),
TO_SIGNED(-57,11),
TO_SIGNED(-103,11),
TO_SIGNED(-150,11),
TO_SIGNED(-195,11),
TO_SIGNED(-240,11),
TO_SIGNED(-284,11),
TO_SIGNED(-327,11),
TO_SIGNED(-369,11),
TO_SIGNED(-409,11),
TO_SIGNED(-448,11),
TO_SIGNED(-485,11),
TO_SIGNED(-519,11),
TO_SIGNED(-552,11),
TO_SIGNED(-583,11),
TO_SIGNED(-611,11),
TO_SIGNED(-637,11),
TO_SIGNED(-661,11),
TO_SIGNED(-682,11),
TO_SIGNED(-700,11),
TO_SIGNED(-716,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-725,11),
TO_SIGNED(-711,11),
TO_SIGNED(-695,11),
TO_SIGNED(-676,11),
TO_SIGNED(-654,11),
TO_SIGNED(-630,11),
TO_SIGNED(-603,11),
TO_SIGNED(-574,11),
TO_SIGNED(-543,11),
TO_SIGNED(-509,11),
TO_SIGNED(-474,11),
TO_SIGNED(-437,11),
TO_SIGNED(-397,11),
TO_SIGNED(-357,11),
TO_SIGNED(-315,11),
TO_SIGNED(-272,11),
TO_SIGNED(-227,11),
TO_SIGNED(-182,11),
TO_SIGNED(-136,11),
TO_SIGNED(-90,11),
TO_SIGNED(-43,11),
TO_SIGNED(4,11),
TO_SIGNED(51,11),
TO_SIGNED(98,11),
TO_SIGNED(144,11),
TO_SIGNED(190,11),
TO_SIGNED(235,11),
TO_SIGNED(279,11),
TO_SIGNED(323,11),
TO_SIGNED(364,11),
TO_SIGNED(405,11),
TO_SIGNED(443,11),
TO_SIGNED(480,11),
TO_SIGNED(516,11),
TO_SIGNED(549,11),
TO_SIGNED(580,11),
TO_SIGNED(608,11),
TO_SIGNED(635,11),
TO_SIGNED(658,11),
TO_SIGNED(680,11),
TO_SIGNED(698,11),
TO_SIGNED(714,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(713,11),
TO_SIGNED(697,11),
TO_SIGNED(678,11),
TO_SIGNED(657,11),
TO_SIGNED(633,11),
TO_SIGNED(606,11),
TO_SIGNED(578,11),
TO_SIGNED(547,11),
TO_SIGNED(513,11),
TO_SIGNED(478,11),
TO_SIGNED(441,11),
TO_SIGNED(402,11),
TO_SIGNED(362,11),
TO_SIGNED(320,11),
TO_SIGNED(276,11),
TO_SIGNED(232,11),
TO_SIGNED(187,11),
TO_SIGNED(141,11),
TO_SIGNED(95,11),
TO_SIGNED(48,11),
TO_SIGNED(1,11),
TO_SIGNED(-46,11),
TO_SIGNED(-93,11),
TO_SIGNED(-139,11),
TO_SIGNED(-185,11),
TO_SIGNED(-230,11),
TO_SIGNED(-275,11),
TO_SIGNED(-318,11),
TO_SIGNED(-360,11),
TO_SIGNED(-400,11),
TO_SIGNED(-439,11),
TO_SIGNED(-476,11),
TO_SIGNED(-512,11),
TO_SIGNED(-545,11),
TO_SIGNED(-576,11),
TO_SIGNED(-605,11),
TO_SIGNED(-632,11),
TO_SIGNED(-656,11),
TO_SIGNED(-677,11),
TO_SIGNED(-696,11),
TO_SIGNED(-712,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-715,11),
TO_SIGNED(-699,11),
TO_SIGNED(-681,11),
TO_SIGNED(-659,11),
TO_SIGNED(-636,11),
TO_SIGNED(-610,11),
TO_SIGNED(-581,11),
TO_SIGNED(-550,11),
TO_SIGNED(-517,11),
TO_SIGNED(-482,11),
TO_SIGNED(-445,11),
TO_SIGNED(-406,11),
TO_SIGNED(-366,11),
TO_SIGNED(-324,11),
TO_SIGNED(-281,11),
TO_SIGNED(-237,11),
TO_SIGNED(-192,11),
TO_SIGNED(-147,11),
TO_SIGNED(-100,11),
TO_SIGNED(-53,11),
TO_SIGNED(-6,11),
TO_SIGNED(41,11),
TO_SIGNED(87,11),
TO_SIGNED(134,11),
TO_SIGNED(180,11),
TO_SIGNED(225,11),
TO_SIGNED(270,11),
TO_SIGNED(313,11),
TO_SIGNED(355,11),
TO_SIGNED(396,11),
TO_SIGNED(435,11),
TO_SIGNED(472,11),
TO_SIGNED(508,11),
TO_SIGNED(541,11),
TO_SIGNED(573,11),
TO_SIGNED(602,11),
TO_SIGNED(629,11),
TO_SIGNED(653,11),
TO_SIGNED(675,11),
TO_SIGNED(694,11),
TO_SIGNED(711,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(729,11),
TO_SIGNED(716,11),
TO_SIGNED(701,11),
TO_SIGNED(683,11),
TO_SIGNED(662,11),
TO_SIGNED(639,11),
TO_SIGNED(613,11),
TO_SIGNED(584,11),
TO_SIGNED(554,11),
TO_SIGNED(521,11),
TO_SIGNED(486,11),
TO_SIGNED(449,11),
TO_SIGNED(411,11),
TO_SIGNED(371,11),
TO_SIGNED(329,11),
TO_SIGNED(286,11),
TO_SIGNED(242,11),
TO_SIGNED(197,11),
TO_SIGNED(152,11),
TO_SIGNED(105,11),
TO_SIGNED(59,11),
TO_SIGNED(12,11),
TO_SIGNED(-35,11),
TO_SIGNED(-82,11),
TO_SIGNED(-129,11),
TO_SIGNED(-175,11),
TO_SIGNED(-220,11),
TO_SIGNED(-265,11),
TO_SIGNED(-308,11),
TO_SIGNED(-350,11),
TO_SIGNED(-391,11),
TO_SIGNED(-430,11),
TO_SIGNED(-468,11),
TO_SIGNED(-504,11),
TO_SIGNED(-538,11),
TO_SIGNED(-569,11),
TO_SIGNED(-599,11),
TO_SIGNED(-626,11),
TO_SIGNED(-651,11),
TO_SIGNED(-673,11),
TO_SIGNED(-692,11),
TO_SIGNED(-709,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-685,11),
TO_SIGNED(-664,11),
TO_SIGNED(-641,11),
TO_SIGNED(-616,11),
TO_SIGNED(-588,11),
TO_SIGNED(-557,11),
TO_SIGNED(-525,11),
TO_SIGNED(-490,11),
TO_SIGNED(-454,11),
TO_SIGNED(-415,11),
TO_SIGNED(-375,11),
TO_SIGNED(-334,11),
TO_SIGNED(-291,11),
TO_SIGNED(-247,11),
TO_SIGNED(-203,11),
TO_SIGNED(-157,11),
TO_SIGNED(-111,11),
TO_SIGNED(-64,11),
TO_SIGNED(-17,11),
TO_SIGNED(30,11),
TO_SIGNED(77,11),
TO_SIGNED(123,11),
TO_SIGNED(169,11),
TO_SIGNED(215,11),
TO_SIGNED(260,11),
TO_SIGNED(303,11),
TO_SIGNED(345,11),
TO_SIGNED(387,11),
TO_SIGNED(426,11),
TO_SIGNED(464,11),
TO_SIGNED(500,11),
TO_SIGNED(534,11),
TO_SIGNED(566,11),
TO_SIGNED(596,11),
TO_SIGNED(623,11),
TO_SIGNED(648,11),
TO_SIGNED(670,11),
TO_SIGNED(690,11),
TO_SIGNED(707,11),
TO_SIGNED(721,11),
TO_SIGNED(733,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(705,11),
TO_SIGNED(687,11),
TO_SIGNED(667,11),
TO_SIGNED(644,11),
TO_SIGNED(619,11),
TO_SIGNED(591,11),
TO_SIGNED(561,11),
TO_SIGNED(529,11),
TO_SIGNED(494,11),
TO_SIGNED(458,11),
TO_SIGNED(420,11),
TO_SIGNED(380,11),
TO_SIGNED(339,11),
TO_SIGNED(296,11),
TO_SIGNED(252,11),
TO_SIGNED(208,11),
TO_SIGNED(162,11),
TO_SIGNED(116,11),
TO_SIGNED(69,11),
TO_SIGNED(22,11),
TO_SIGNED(-25,11),
TO_SIGNED(-71,11),
TO_SIGNED(-118,11),
TO_SIGNED(-164,11),
TO_SIGNED(-210,11),
TO_SIGNED(-255,11),
TO_SIGNED(-298,11),
TO_SIGNED(-341,11),
TO_SIGNED(-382,11),
TO_SIGNED(-422,11),
TO_SIGNED(-460,11),
TO_SIGNED(-496,11),
TO_SIGNED(-530,11),
TO_SIGNED(-562,11),
TO_SIGNED(-592,11),
TO_SIGNED(-620,11),
TO_SIGNED(-645,11),
TO_SIGNED(-668,11),
TO_SIGNED(-688,11),
TO_SIGNED(-705,11),
TO_SIGNED(-720,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-721,11),
TO_SIGNED(-706,11),
TO_SIGNED(-689,11),
TO_SIGNED(-669,11),
TO_SIGNED(-647,11),
TO_SIGNED(-622,11),
TO_SIGNED(-594,11),
TO_SIGNED(-564,11),
TO_SIGNED(-532,11),
TO_SIGNED(-498,11),
TO_SIGNED(-462,11),
TO_SIGNED(-424,11),
TO_SIGNED(-385,11),
TO_SIGNED(-344,11),
TO_SIGNED(-301,11),
TO_SIGNED(-258,11),
TO_SIGNED(-213,11),
TO_SIGNED(-167,11),
TO_SIGNED(-121,11),
TO_SIGNED(-75,11),
TO_SIGNED(-28,11),
TO_SIGNED(19,11),
TO_SIGNED(66,11),
TO_SIGNED(113,11),
TO_SIGNED(159,11),
TO_SIGNED(205,11),
TO_SIGNED(249,11),
TO_SIGNED(293,11),
TO_SIGNED(336,11),
TO_SIGNED(377,11),
TO_SIGNED(417,11),
TO_SIGNED(455,11),
TO_SIGNED(492,11),
TO_SIGNED(526,11),
TO_SIGNED(559,11),
TO_SIGNED(589,11),
TO_SIGNED(617,11),
TO_SIGNED(642,11),
TO_SIGNED(665,11),
TO_SIGNED(686,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(708,11),
TO_SIGNED(691,11),
TO_SIGNED(672,11),
TO_SIGNED(650,11),
TO_SIGNED(625,11),
TO_SIGNED(598,11),
TO_SIGNED(568,11),
TO_SIGNED(536,11),
TO_SIGNED(502,11),
TO_SIGNED(466,11),
TO_SIGNED(429,11),
TO_SIGNED(389,11),
TO_SIGNED(348,11),
TO_SIGNED(306,11),
TO_SIGNED(263,11),
TO_SIGNED(218,11),
TO_SIGNED(173,11),
TO_SIGNED(127,11),
TO_SIGNED(80,11),
TO_SIGNED(33,11),
TO_SIGNED(-14,11),
TO_SIGNED(-61,11),
TO_SIGNED(-108,11),
TO_SIGNED(-154,11),
TO_SIGNED(-200,11),
TO_SIGNED(-244,11),
TO_SIGNED(-288,11),
TO_SIGNED(-331,11),
TO_SIGNED(-373,11),
TO_SIGNED(-413,11),
TO_SIGNED(-451,11),
TO_SIGNED(-488,11),
TO_SIGNED(-523,11),
TO_SIGNED(-555,11),
TO_SIGNED(-586,11),
TO_SIGNED(-614,11),
TO_SIGNED(-640,11),
TO_SIGNED(-663,11),
TO_SIGNED(-684,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-729,11),
TO_SIGNED(-739,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-710,11),
TO_SIGNED(-693,11),
TO_SIGNED(-674,11),
TO_SIGNED(-652,11),
TO_SIGNED(-628,11),
TO_SIGNED(-601,11),
TO_SIGNED(-571,11),
TO_SIGNED(-540,11),
TO_SIGNED(-506,11),
TO_SIGNED(-471,11),
TO_SIGNED(-433,11),
TO_SIGNED(-394,11),
TO_SIGNED(-353,11),
TO_SIGNED(-311,11),
TO_SIGNED(-268,11),
TO_SIGNED(-223,11),
TO_SIGNED(-178,11),
TO_SIGNED(-132,11),
TO_SIGNED(-85,11),
TO_SIGNED(-38,11),
TO_SIGNED(9,11),
TO_SIGNED(56,11),
TO_SIGNED(102,11),
TO_SIGNED(149,11),
TO_SIGNED(194,11),
TO_SIGNED(239,11),
TO_SIGNED(283,11),
TO_SIGNED(326,11),
TO_SIGNED(368,11),
TO_SIGNED(408,11),
TO_SIGNED(447,11),
TO_SIGNED(484,11),
TO_SIGNED(519,11),
TO_SIGNED(552,11),
TO_SIGNED(582,11),
TO_SIGNED(611,11),
TO_SIGNED(637,11),
TO_SIGNED(660,11),
TO_SIGNED(681,11),
TO_SIGNED(700,11),
TO_SIGNED(715,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(736,11),
TO_SIGNED(725,11),
TO_SIGNED(712,11),
TO_SIGNED(695,11),
TO_SIGNED(676,11),
TO_SIGNED(655,11),
TO_SIGNED(631,11),
TO_SIGNED(604,11),
TO_SIGNED(575,11),
TO_SIGNED(544,11),
TO_SIGNED(510,11),
TO_SIGNED(475,11),
TO_SIGNED(437,11),
TO_SIGNED(398,11),
TO_SIGNED(358,11),
TO_SIGNED(316,11),
TO_SIGNED(273,11),
TO_SIGNED(228,11),
TO_SIGNED(183,11),
TO_SIGNED(137,11),
TO_SIGNED(91,11),
TO_SIGNED(44,11),
TO_SIGNED(-3,11),
TO_SIGNED(-50,11),
TO_SIGNED(-97,11),
TO_SIGNED(-143,11),
TO_SIGNED(-189,11),
TO_SIGNED(-234,11),
TO_SIGNED(-278,11),
TO_SIGNED(-322,11),
TO_SIGNED(-363,11),
TO_SIGNED(-404,11),
TO_SIGNED(-443,11),
TO_SIGNED(-480,11),
TO_SIGNED(-515,11),
TO_SIGNED(-548,11),
TO_SIGNED(-579,11),
TO_SIGNED(-608,11),
TO_SIGNED(-634,11),
TO_SIGNED(-658,11),
TO_SIGNED(-679,11),
TO_SIGNED(-698,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-679,11),
TO_SIGNED(-657,11),
TO_SIGNED(-633,11),
TO_SIGNED(-607,11),
TO_SIGNED(-578,11),
TO_SIGNED(-547,11),
TO_SIGNED(-514,11),
TO_SIGNED(-479,11),
TO_SIGNED(-442,11),
TO_SIGNED(-403,11),
TO_SIGNED(-362,11),
TO_SIGNED(-321,11),
TO_SIGNED(-277,11),
TO_SIGNED(-233,11),
TO_SIGNED(-188,11),
TO_SIGNED(-142,11),
TO_SIGNED(-96,11),
TO_SIGNED(-49,11),
TO_SIGNED(-2,11),
TO_SIGNED(45,11),
TO_SIGNED(92,11),
TO_SIGNED(138,11),
TO_SIGNED(184,11),
TO_SIGNED(229,11),
TO_SIGNED(274,11),
TO_SIGNED(317,11),
TO_SIGNED(359,11),
TO_SIGNED(399,11),
TO_SIGNED(438,11),
TO_SIGNED(476,11),
TO_SIGNED(511,11),
TO_SIGNED(544,11),
TO_SIGNED(576,11),
TO_SIGNED(605,11),
TO_SIGNED(631,11),
TO_SIGNED(655,11),
TO_SIGNED(677,11),
TO_SIGNED(696,11),
TO_SIGNED(712,11),
TO_SIGNED(725,11),
TO_SIGNED(736,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(715,11),
TO_SIGNED(699,11),
TO_SIGNED(681,11),
TO_SIGNED(660,11),
TO_SIGNED(636,11),
TO_SIGNED(610,11),
TO_SIGNED(582,11),
TO_SIGNED(551,11),
TO_SIGNED(518,11),
TO_SIGNED(483,11),
TO_SIGNED(446,11),
TO_SIGNED(407,11),
TO_SIGNED(367,11),
TO_SIGNED(325,11),
TO_SIGNED(282,11),
TO_SIGNED(238,11),
TO_SIGNED(193,11),
TO_SIGNED(148,11),
TO_SIGNED(101,11),
TO_SIGNED(54,11),
TO_SIGNED(7,11),
TO_SIGNED(-40,11),
TO_SIGNED(-86,11),
TO_SIGNED(-133,11),
TO_SIGNED(-179,11),
TO_SIGNED(-224,11),
TO_SIGNED(-269,11),
TO_SIGNED(-312,11),
TO_SIGNED(-354,11),
TO_SIGNED(-395,11),
TO_SIGNED(-434,11),
TO_SIGNED(-471,11),
TO_SIGNED(-507,11),
TO_SIGNED(-541,11),
TO_SIGNED(-572,11),
TO_SIGNED(-601,11),
TO_SIGNED(-628,11),
TO_SIGNED(-653,11),
TO_SIGNED(-675,11),
TO_SIGNED(-694,11),
TO_SIGNED(-710,11),
TO_SIGNED(-724,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-701,11),
TO_SIGNED(-683,11),
TO_SIGNED(-662,11),
TO_SIGNED(-639,11),
TO_SIGNED(-613,11),
TO_SIGNED(-585,11),
TO_SIGNED(-554,11),
TO_SIGNED(-522,11),
TO_SIGNED(-487,11),
TO_SIGNED(-450,11),
TO_SIGNED(-412,11),
TO_SIGNED(-372,11),
TO_SIGNED(-330,11),
TO_SIGNED(-287,11),
TO_SIGNED(-243,11),
TO_SIGNED(-198,11),
TO_SIGNED(-153,11),
TO_SIGNED(-106,11),
TO_SIGNED(-60,11),
TO_SIGNED(-13,11),
TO_SIGNED(34,11),
TO_SIGNED(81,11),
TO_SIGNED(128,11),
TO_SIGNED(174,11),
TO_SIGNED(219,11),
TO_SIGNED(264,11),
TO_SIGNED(307,11),
TO_SIGNED(349,11),
TO_SIGNED(390,11),
TO_SIGNED(430,11),
TO_SIGNED(467,11),
TO_SIGNED(503,11),
TO_SIGNED(537,11),
TO_SIGNED(569,11),
TO_SIGNED(598,11),
TO_SIGNED(625,11),
TO_SIGNED(650,11),
TO_SIGNED(672,11),
TO_SIGNED(692,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(730,11),
TO_SIGNED(718,11),
TO_SIGNED(703,11),
TO_SIGNED(685,11),
TO_SIGNED(665,11),
TO_SIGNED(642,11),
TO_SIGNED(616,11),
TO_SIGNED(588,11),
TO_SIGNED(558,11),
TO_SIGNED(526,11),
TO_SIGNED(491,11),
TO_SIGNED(455,11),
TO_SIGNED(416,11),
TO_SIGNED(376,11),
TO_SIGNED(335,11),
TO_SIGNED(292,11),
TO_SIGNED(248,11),
TO_SIGNED(204,11),
TO_SIGNED(158,11),
TO_SIGNED(112,11),
TO_SIGNED(65,11),
TO_SIGNED(18,11),
TO_SIGNED(-29,11),
TO_SIGNED(-76,11),
TO_SIGNED(-122,11),
TO_SIGNED(-168,11),
TO_SIGNED(-214,11),
TO_SIGNED(-259,11),
TO_SIGNED(-302,11),
TO_SIGNED(-345,11),
TO_SIGNED(-386,11),
TO_SIGNED(-425,11),
TO_SIGNED(-463,11),
TO_SIGNED(-499,11),
TO_SIGNED(-533,11),
TO_SIGNED(-565,11),
TO_SIGNED(-595,11),
TO_SIGNED(-622,11),
TO_SIGNED(-647,11),
TO_SIGNED(-670,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-721,11),
TO_SIGNED(-733,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-720,11),
TO_SIGNED(-705,11),
TO_SIGNED(-688,11),
TO_SIGNED(-667,11),
TO_SIGNED(-645,11),
TO_SIGNED(-619,11),
TO_SIGNED(-592,11),
TO_SIGNED(-562,11),
TO_SIGNED(-529,11),
TO_SIGNED(-495,11),
TO_SIGNED(-459,11),
TO_SIGNED(-421,11),
TO_SIGNED(-381,11),
TO_SIGNED(-340,11),
TO_SIGNED(-297,11),
TO_SIGNED(-254,11),
TO_SIGNED(-209,11),
TO_SIGNED(-163,11),
TO_SIGNED(-117,11),
TO_SIGNED(-70,11),
TO_SIGNED(-24,11),
TO_SIGNED(24,11),
TO_SIGNED(70,11),
TO_SIGNED(117,11),
TO_SIGNED(163,11),
TO_SIGNED(209,11),
TO_SIGNED(254,11),
TO_SIGNED(297,11),
TO_SIGNED(340,11),
TO_SIGNED(381,11),
TO_SIGNED(421,11),
TO_SIGNED(459,11),
TO_SIGNED(495,11),
TO_SIGNED(529,11),
TO_SIGNED(562,11),
TO_SIGNED(592,11),
TO_SIGNED(619,11),
TO_SIGNED(645,11),
TO_SIGNED(667,11),
TO_SIGNED(688,11),
TO_SIGNED(705,11),
TO_SIGNED(720,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(733,11),
TO_SIGNED(721,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(670,11),
TO_SIGNED(647,11),
TO_SIGNED(622,11),
TO_SIGNED(595,11),
TO_SIGNED(565,11),
TO_SIGNED(533,11),
TO_SIGNED(499,11),
TO_SIGNED(463,11),
TO_SIGNED(425,11),
TO_SIGNED(386,11),
TO_SIGNED(345,11),
TO_SIGNED(302,11),
TO_SIGNED(259,11),
TO_SIGNED(214,11),
TO_SIGNED(168,11),
TO_SIGNED(122,11),
TO_SIGNED(76,11),
TO_SIGNED(29,11),
TO_SIGNED(-18,11),
TO_SIGNED(-65,11),
TO_SIGNED(-112,11),
TO_SIGNED(-158,11),
TO_SIGNED(-204,11),
TO_SIGNED(-248,11),
TO_SIGNED(-292,11),
TO_SIGNED(-335,11),
TO_SIGNED(-376,11),
TO_SIGNED(-416,11),
TO_SIGNED(-455,11),
TO_SIGNED(-491,11),
TO_SIGNED(-526,11),
TO_SIGNED(-558,11),
TO_SIGNED(-588,11),
TO_SIGNED(-616,11),
TO_SIGNED(-642,11),
TO_SIGNED(-665,11),
TO_SIGNED(-685,11),
TO_SIGNED(-703,11),
TO_SIGNED(-718,11),
TO_SIGNED(-730,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-692,11),
TO_SIGNED(-672,11),
TO_SIGNED(-650,11),
TO_SIGNED(-625,11),
TO_SIGNED(-598,11),
TO_SIGNED(-569,11),
TO_SIGNED(-537,11),
TO_SIGNED(-503,11),
TO_SIGNED(-467,11),
TO_SIGNED(-430,11),
TO_SIGNED(-390,11),
TO_SIGNED(-349,11),
TO_SIGNED(-307,11),
TO_SIGNED(-264,11),
TO_SIGNED(-219,11),
TO_SIGNED(-174,11),
TO_SIGNED(-128,11),
TO_SIGNED(-81,11),
TO_SIGNED(-34,11),
TO_SIGNED(13,11),
TO_SIGNED(60,11),
TO_SIGNED(106,11),
TO_SIGNED(153,11),
TO_SIGNED(198,11),
TO_SIGNED(243,11),
TO_SIGNED(287,11),
TO_SIGNED(330,11),
TO_SIGNED(372,11),
TO_SIGNED(412,11),
TO_SIGNED(450,11),
TO_SIGNED(487,11),
TO_SIGNED(522,11),
TO_SIGNED(554,11),
TO_SIGNED(585,11),
TO_SIGNED(613,11),
TO_SIGNED(639,11),
TO_SIGNED(662,11),
TO_SIGNED(683,11),
TO_SIGNED(701,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(724,11),
TO_SIGNED(710,11),
TO_SIGNED(694,11),
TO_SIGNED(675,11),
TO_SIGNED(653,11),
TO_SIGNED(628,11),
TO_SIGNED(601,11),
TO_SIGNED(572,11),
TO_SIGNED(541,11),
TO_SIGNED(507,11),
TO_SIGNED(471,11),
TO_SIGNED(434,11),
TO_SIGNED(395,11),
TO_SIGNED(354,11),
TO_SIGNED(312,11),
TO_SIGNED(269,11),
TO_SIGNED(224,11),
TO_SIGNED(179,11),
TO_SIGNED(133,11),
TO_SIGNED(86,11),
TO_SIGNED(40,11),
TO_SIGNED(-7,11),
TO_SIGNED(-54,11),
TO_SIGNED(-101,11),
TO_SIGNED(-148,11),
TO_SIGNED(-193,11),
TO_SIGNED(-238,11),
TO_SIGNED(-282,11),
TO_SIGNED(-325,11),
TO_SIGNED(-367,11),
TO_SIGNED(-407,11),
TO_SIGNED(-446,11),
TO_SIGNED(-483,11),
TO_SIGNED(-518,11),
TO_SIGNED(-551,11),
TO_SIGNED(-582,11),
TO_SIGNED(-610,11),
TO_SIGNED(-636,11),
TO_SIGNED(-660,11),
TO_SIGNED(-681,11),
TO_SIGNED(-699,11),
TO_SIGNED(-715,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-736,11),
TO_SIGNED(-725,11),
TO_SIGNED(-712,11),
TO_SIGNED(-696,11),
TO_SIGNED(-677,11),
TO_SIGNED(-655,11),
TO_SIGNED(-631,11),
TO_SIGNED(-605,11),
TO_SIGNED(-576,11),
TO_SIGNED(-544,11),
TO_SIGNED(-511,11),
TO_SIGNED(-476,11),
TO_SIGNED(-438,11),
TO_SIGNED(-399,11),
TO_SIGNED(-359,11),
TO_SIGNED(-317,11),
TO_SIGNED(-274,11),
TO_SIGNED(-229,11),
TO_SIGNED(-184,11),
TO_SIGNED(-138,11),
TO_SIGNED(-92,11),
TO_SIGNED(-45,11),
TO_SIGNED(2,11),
TO_SIGNED(49,11),
TO_SIGNED(96,11),
TO_SIGNED(142,11),
TO_SIGNED(188,11),
TO_SIGNED(233,11),
TO_SIGNED(277,11),
TO_SIGNED(321,11),
TO_SIGNED(362,11),
TO_SIGNED(403,11),
TO_SIGNED(442,11),
TO_SIGNED(479,11),
TO_SIGNED(514,11),
TO_SIGNED(547,11),
TO_SIGNED(578,11),
TO_SIGNED(607,11),
TO_SIGNED(633,11),
TO_SIGNED(657,11),
TO_SIGNED(679,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(698,11),
TO_SIGNED(679,11),
TO_SIGNED(658,11),
TO_SIGNED(634,11),
TO_SIGNED(608,11),
TO_SIGNED(579,11),
TO_SIGNED(548,11),
TO_SIGNED(515,11),
TO_SIGNED(480,11),
TO_SIGNED(443,11),
TO_SIGNED(404,11),
TO_SIGNED(363,11),
TO_SIGNED(322,11),
TO_SIGNED(278,11),
TO_SIGNED(234,11),
TO_SIGNED(189,11),
TO_SIGNED(143,11),
TO_SIGNED(97,11),
TO_SIGNED(50,11),
TO_SIGNED(3,11),
TO_SIGNED(-44,11),
TO_SIGNED(-91,11),
TO_SIGNED(-137,11),
TO_SIGNED(-183,11),
TO_SIGNED(-228,11),
TO_SIGNED(-273,11),
TO_SIGNED(-316,11),
TO_SIGNED(-358,11),
TO_SIGNED(-398,11),
TO_SIGNED(-437,11),
TO_SIGNED(-475,11),
TO_SIGNED(-510,11),
TO_SIGNED(-544,11),
TO_SIGNED(-575,11),
TO_SIGNED(-604,11),
TO_SIGNED(-631,11),
TO_SIGNED(-655,11),
TO_SIGNED(-676,11),
TO_SIGNED(-695,11),
TO_SIGNED(-712,11),
TO_SIGNED(-725,11),
TO_SIGNED(-736,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-715,11),
TO_SIGNED(-700,11),
TO_SIGNED(-681,11),
TO_SIGNED(-660,11),
TO_SIGNED(-637,11),
TO_SIGNED(-611,11),
TO_SIGNED(-582,11),
TO_SIGNED(-552,11),
TO_SIGNED(-519,11),
TO_SIGNED(-484,11),
TO_SIGNED(-447,11),
TO_SIGNED(-408,11),
TO_SIGNED(-368,11),
TO_SIGNED(-326,11),
TO_SIGNED(-283,11),
TO_SIGNED(-239,11),
TO_SIGNED(-194,11),
TO_SIGNED(-149,11),
TO_SIGNED(-102,11),
TO_SIGNED(-56,11),
TO_SIGNED(-9,11),
TO_SIGNED(38,11),
TO_SIGNED(85,11),
TO_SIGNED(132,11),
TO_SIGNED(178,11),
TO_SIGNED(223,11),
TO_SIGNED(268,11),
TO_SIGNED(311,11),
TO_SIGNED(353,11),
TO_SIGNED(394,11),
TO_SIGNED(433,11),
TO_SIGNED(471,11),
TO_SIGNED(506,11),
TO_SIGNED(540,11),
TO_SIGNED(571,11),
TO_SIGNED(601,11),
TO_SIGNED(628,11),
TO_SIGNED(652,11),
TO_SIGNED(674,11),
TO_SIGNED(693,11),
TO_SIGNED(710,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(739,11),
TO_SIGNED(729,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(684,11),
TO_SIGNED(663,11),
TO_SIGNED(640,11),
TO_SIGNED(614,11),
TO_SIGNED(586,11),
TO_SIGNED(555,11),
TO_SIGNED(523,11),
TO_SIGNED(488,11),
TO_SIGNED(451,11),
TO_SIGNED(413,11),
TO_SIGNED(373,11),
TO_SIGNED(331,11),
TO_SIGNED(288,11),
TO_SIGNED(244,11),
TO_SIGNED(200,11),
TO_SIGNED(154,11),
TO_SIGNED(108,11),
TO_SIGNED(61,11),
TO_SIGNED(14,11),
TO_SIGNED(-33,11),
TO_SIGNED(-80,11),
TO_SIGNED(-127,11),
TO_SIGNED(-173,11),
TO_SIGNED(-218,11),
TO_SIGNED(-263,11),
TO_SIGNED(-306,11),
TO_SIGNED(-348,11),
TO_SIGNED(-389,11),
TO_SIGNED(-429,11),
TO_SIGNED(-466,11),
TO_SIGNED(-502,11),
TO_SIGNED(-536,11),
TO_SIGNED(-568,11),
TO_SIGNED(-598,11),
TO_SIGNED(-625,11),
TO_SIGNED(-650,11),
TO_SIGNED(-672,11),
TO_SIGNED(-691,11),
TO_SIGNED(-708,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-686,11),
TO_SIGNED(-665,11),
TO_SIGNED(-642,11),
TO_SIGNED(-617,11),
TO_SIGNED(-589,11),
TO_SIGNED(-559,11),
TO_SIGNED(-526,11),
TO_SIGNED(-492,11),
TO_SIGNED(-455,11),
TO_SIGNED(-417,11),
TO_SIGNED(-377,11),
TO_SIGNED(-336,11),
TO_SIGNED(-293,11),
TO_SIGNED(-249,11),
TO_SIGNED(-205,11),
TO_SIGNED(-159,11),
TO_SIGNED(-113,11),
TO_SIGNED(-66,11),
TO_SIGNED(-19,11),
TO_SIGNED(28,11),
TO_SIGNED(75,11),
TO_SIGNED(121,11),
TO_SIGNED(167,11),
TO_SIGNED(213,11),
TO_SIGNED(258,11),
TO_SIGNED(301,11),
TO_SIGNED(344,11),
TO_SIGNED(385,11),
TO_SIGNED(424,11),
TO_SIGNED(462,11),
TO_SIGNED(498,11),
TO_SIGNED(532,11),
TO_SIGNED(564,11),
TO_SIGNED(594,11),
TO_SIGNED(622,11),
TO_SIGNED(647,11),
TO_SIGNED(669,11),
TO_SIGNED(689,11),
TO_SIGNED(706,11),
TO_SIGNED(721,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(720,11),
TO_SIGNED(705,11),
TO_SIGNED(688,11),
TO_SIGNED(668,11),
TO_SIGNED(645,11),
TO_SIGNED(620,11),
TO_SIGNED(592,11),
TO_SIGNED(562,11),
TO_SIGNED(530,11),
TO_SIGNED(496,11),
TO_SIGNED(460,11),
TO_SIGNED(422,11),
TO_SIGNED(382,11),
TO_SIGNED(341,11),
TO_SIGNED(298,11),
TO_SIGNED(255,11),
TO_SIGNED(210,11),
TO_SIGNED(164,11),
TO_SIGNED(118,11),
TO_SIGNED(71,11),
TO_SIGNED(25,11),
TO_SIGNED(-22,11),
TO_SIGNED(-69,11),
TO_SIGNED(-116,11),
TO_SIGNED(-162,11),
TO_SIGNED(-208,11),
TO_SIGNED(-252,11),
TO_SIGNED(-296,11),
TO_SIGNED(-339,11),
TO_SIGNED(-380,11),
TO_SIGNED(-420,11),
TO_SIGNED(-458,11),
TO_SIGNED(-494,11),
TO_SIGNED(-529,11),
TO_SIGNED(-561,11),
TO_SIGNED(-591,11),
TO_SIGNED(-619,11),
TO_SIGNED(-644,11),
TO_SIGNED(-667,11),
TO_SIGNED(-687,11),
TO_SIGNED(-705,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-733,11),
TO_SIGNED(-721,11),
TO_SIGNED(-707,11),
TO_SIGNED(-690,11),
TO_SIGNED(-670,11),
TO_SIGNED(-648,11),
TO_SIGNED(-623,11),
TO_SIGNED(-596,11),
TO_SIGNED(-566,11),
TO_SIGNED(-534,11),
TO_SIGNED(-500,11),
TO_SIGNED(-464,11),
TO_SIGNED(-426,11),
TO_SIGNED(-387,11),
TO_SIGNED(-345,11),
TO_SIGNED(-303,11),
TO_SIGNED(-260,11),
TO_SIGNED(-215,11),
TO_SIGNED(-169,11),
TO_SIGNED(-123,11),
TO_SIGNED(-77,11),
TO_SIGNED(-30,11),
TO_SIGNED(17,11),
TO_SIGNED(64,11),
TO_SIGNED(111,11),
TO_SIGNED(157,11),
TO_SIGNED(203,11),
TO_SIGNED(247,11),
TO_SIGNED(291,11),
TO_SIGNED(334,11),
TO_SIGNED(375,11),
TO_SIGNED(415,11),
TO_SIGNED(454,11),
TO_SIGNED(490,11),
TO_SIGNED(525,11),
TO_SIGNED(557,11),
TO_SIGNED(588,11),
TO_SIGNED(616,11),
TO_SIGNED(641,11),
TO_SIGNED(664,11),
TO_SIGNED(685,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(709,11),
TO_SIGNED(692,11),
TO_SIGNED(673,11),
TO_SIGNED(651,11),
TO_SIGNED(626,11),
TO_SIGNED(599,11),
TO_SIGNED(569,11),
TO_SIGNED(538,11),
TO_SIGNED(504,11),
TO_SIGNED(468,11),
TO_SIGNED(430,11),
TO_SIGNED(391,11),
TO_SIGNED(350,11),
TO_SIGNED(308,11),
TO_SIGNED(265,11),
TO_SIGNED(220,11),
TO_SIGNED(175,11),
TO_SIGNED(129,11),
TO_SIGNED(82,11),
TO_SIGNED(35,11),
TO_SIGNED(-12,11),
TO_SIGNED(-59,11),
TO_SIGNED(-105,11),
TO_SIGNED(-152,11),
TO_SIGNED(-197,11),
TO_SIGNED(-242,11),
TO_SIGNED(-286,11),
TO_SIGNED(-329,11),
TO_SIGNED(-371,11),
TO_SIGNED(-411,11),
TO_SIGNED(-449,11),
TO_SIGNED(-486,11),
TO_SIGNED(-521,11),
TO_SIGNED(-554,11),
TO_SIGNED(-584,11),
TO_SIGNED(-613,11),
TO_SIGNED(-639,11),
TO_SIGNED(-662,11),
TO_SIGNED(-683,11),
TO_SIGNED(-701,11),
TO_SIGNED(-716,11),
TO_SIGNED(-729,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-711,11),
TO_SIGNED(-694,11),
TO_SIGNED(-675,11),
TO_SIGNED(-653,11),
TO_SIGNED(-629,11),
TO_SIGNED(-602,11),
TO_SIGNED(-573,11),
TO_SIGNED(-541,11),
TO_SIGNED(-508,11),
TO_SIGNED(-472,11),
TO_SIGNED(-435,11),
TO_SIGNED(-396,11),
TO_SIGNED(-355,11),
TO_SIGNED(-313,11),
TO_SIGNED(-270,11),
TO_SIGNED(-225,11),
TO_SIGNED(-180,11),
TO_SIGNED(-134,11),
TO_SIGNED(-87,11),
TO_SIGNED(-41,11),
TO_SIGNED(6,11),
TO_SIGNED(53,11),
TO_SIGNED(100,11),
TO_SIGNED(147,11),
TO_SIGNED(192,11),
TO_SIGNED(237,11),
TO_SIGNED(281,11),
TO_SIGNED(324,11),
TO_SIGNED(366,11),
TO_SIGNED(406,11),
TO_SIGNED(445,11),
TO_SIGNED(482,11),
TO_SIGNED(517,11),
TO_SIGNED(550,11),
TO_SIGNED(581,11),
TO_SIGNED(610,11),
TO_SIGNED(636,11),
TO_SIGNED(659,11),
TO_SIGNED(681,11),
TO_SIGNED(699,11),
TO_SIGNED(715,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(712,11),
TO_SIGNED(696,11),
TO_SIGNED(677,11),
TO_SIGNED(656,11),
TO_SIGNED(632,11),
TO_SIGNED(605,11),
TO_SIGNED(576,11),
TO_SIGNED(545,11),
TO_SIGNED(512,11),
TO_SIGNED(476,11),
TO_SIGNED(439,11),
TO_SIGNED(400,11),
TO_SIGNED(360,11),
TO_SIGNED(318,11),
TO_SIGNED(275,11),
TO_SIGNED(230,11),
TO_SIGNED(185,11),
TO_SIGNED(139,11),
TO_SIGNED(93,11),
TO_SIGNED(46,11),
TO_SIGNED(-1,11),
TO_SIGNED(-48,11),
TO_SIGNED(-95,11),
TO_SIGNED(-141,11),
TO_SIGNED(-187,11),
TO_SIGNED(-232,11),
TO_SIGNED(-276,11),
TO_SIGNED(-320,11),
TO_SIGNED(-362,11),
TO_SIGNED(-402,11),
TO_SIGNED(-441,11),
TO_SIGNED(-478,11),
TO_SIGNED(-513,11),
TO_SIGNED(-547,11),
TO_SIGNED(-578,11),
TO_SIGNED(-606,11),
TO_SIGNED(-633,11),
TO_SIGNED(-657,11),
TO_SIGNED(-678,11),
TO_SIGNED(-697,11),
TO_SIGNED(-713,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-714,11),
TO_SIGNED(-698,11),
TO_SIGNED(-680,11),
TO_SIGNED(-658,11),
TO_SIGNED(-635,11),
TO_SIGNED(-608,11),
TO_SIGNED(-580,11),
TO_SIGNED(-549,11),
TO_SIGNED(-516,11),
TO_SIGNED(-480,11),
TO_SIGNED(-443,11),
TO_SIGNED(-405,11),
TO_SIGNED(-364,11),
TO_SIGNED(-323,11),
TO_SIGNED(-279,11),
TO_SIGNED(-235,11),
TO_SIGNED(-190,11),
TO_SIGNED(-144,11),
TO_SIGNED(-98,11),
TO_SIGNED(-51,11),
TO_SIGNED(-4,11),
TO_SIGNED(43,11),
TO_SIGNED(90,11),
TO_SIGNED(136,11),
TO_SIGNED(182,11),
TO_SIGNED(227,11),
TO_SIGNED(272,11),
TO_SIGNED(315,11),
TO_SIGNED(357,11),
TO_SIGNED(397,11),
TO_SIGNED(437,11),
TO_SIGNED(474,11),
TO_SIGNED(509,11),
TO_SIGNED(543,11),
TO_SIGNED(574,11),
TO_SIGNED(603,11),
TO_SIGNED(630,11),
TO_SIGNED(654,11),
TO_SIGNED(676,11),
TO_SIGNED(695,11),
TO_SIGNED(711,11),
TO_SIGNED(725,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(716,11),
TO_SIGNED(700,11),
TO_SIGNED(682,11),
TO_SIGNED(661,11),
TO_SIGNED(637,11),
TO_SIGNED(611,11),
TO_SIGNED(583,11),
TO_SIGNED(552,11),
TO_SIGNED(519,11),
TO_SIGNED(485,11),
TO_SIGNED(448,11),
TO_SIGNED(409,11),
TO_SIGNED(369,11),
TO_SIGNED(327,11),
TO_SIGNED(284,11),
TO_SIGNED(240,11),
TO_SIGNED(195,11),
TO_SIGNED(150,11),
TO_SIGNED(103,11),
TO_SIGNED(57,11),
TO_SIGNED(10,11),
TO_SIGNED(-37,11),
TO_SIGNED(-84,11),
TO_SIGNED(-131,11),
TO_SIGNED(-177,11),
TO_SIGNED(-222,11),
TO_SIGNED(-267,11),
TO_SIGNED(-310,11),
TO_SIGNED(-352,11),
TO_SIGNED(-393,11),
TO_SIGNED(-432,11),
TO_SIGNED(-470,11),
TO_SIGNED(-505,11),
TO_SIGNED(-539,11),
TO_SIGNED(-571,11),
TO_SIGNED(-600,11),
TO_SIGNED(-627,11),
TO_SIGNED(-652,11),
TO_SIGNED(-674,11),
TO_SIGNED(-693,11),
TO_SIGNED(-710,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-702,11),
TO_SIGNED(-684,11),
TO_SIGNED(-663,11),
TO_SIGNED(-640,11),
TO_SIGNED(-615,11),
TO_SIGNED(-586,11),
TO_SIGNED(-556,11),
TO_SIGNED(-523,11),
TO_SIGNED(-489,11),
TO_SIGNED(-452,11),
TO_SIGNED(-414,11),
TO_SIGNED(-374,11),
TO_SIGNED(-332,11),
TO_SIGNED(-289,11),
TO_SIGNED(-245,11),
TO_SIGNED(-201,11),
TO_SIGNED(-155,11),
TO_SIGNED(-109,11),
TO_SIGNED(-62,11),
TO_SIGNED(-15,11),
TO_SIGNED(32,11),
TO_SIGNED(79,11),
TO_SIGNED(125,11),
TO_SIGNED(172,11),
TO_SIGNED(217,11),
TO_SIGNED(262,11),
TO_SIGNED(305,11),
TO_SIGNED(347,11),
TO_SIGNED(388,11),
TO_SIGNED(428,11),
TO_SIGNED(466,11),
TO_SIGNED(501,11),
TO_SIGNED(535,11),
TO_SIGNED(567,11),
TO_SIGNED(597,11),
TO_SIGNED(624,11),
TO_SIGNED(649,11),
TO_SIGNED(671,11),
TO_SIGNED(691,11),
TO_SIGNED(708,11),
TO_SIGNED(722,11),
TO_SIGNED(733,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(704,11),
TO_SIGNED(686,11),
TO_SIGNED(666,11),
TO_SIGNED(643,11),
TO_SIGNED(618,11),
TO_SIGNED(590,11),
TO_SIGNED(559,11),
TO_SIGNED(527,11),
TO_SIGNED(493,11),
TO_SIGNED(456,11),
TO_SIGNED(418,11),
TO_SIGNED(378,11),
TO_SIGNED(337,11),
TO_SIGNED(294,11),
TO_SIGNED(250,11),
TO_SIGNED(206,11),
TO_SIGNED(160,11),
TO_SIGNED(114,11),
TO_SIGNED(67,11),
TO_SIGNED(20,11),
TO_SIGNED(-27,11),
TO_SIGNED(-74,11),
TO_SIGNED(-120,11),
TO_SIGNED(-166,11),
TO_SIGNED(-212,11),
TO_SIGNED(-257,11),
TO_SIGNED(-300,11),
TO_SIGNED(-343,11),
TO_SIGNED(-384,11),
TO_SIGNED(-423,11),
TO_SIGNED(-461,11),
TO_SIGNED(-497,11),
TO_SIGNED(-532,11),
TO_SIGNED(-564,11),
TO_SIGNED(-594,11),
TO_SIGNED(-621,11),
TO_SIGNED(-646,11),
TO_SIGNED(-669,11),
TO_SIGNED(-689,11),
TO_SIGNED(-706,11),
TO_SIGNED(-721,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-720,11),
TO_SIGNED(-706,11),
TO_SIGNED(-688,11),
TO_SIGNED(-668,11),
TO_SIGNED(-646,11),
TO_SIGNED(-621,11),
TO_SIGNED(-593,11),
TO_SIGNED(-563,11),
TO_SIGNED(-531,11),
TO_SIGNED(-497,11),
TO_SIGNED(-460,11),
TO_SIGNED(-422,11),
TO_SIGNED(-383,11),
TO_SIGNED(-342,11),
TO_SIGNED(-299,11),
TO_SIGNED(-256,11),
TO_SIGNED(-211,11),
TO_SIGNED(-165,11),
TO_SIGNED(-119,11),
TO_SIGNED(-73,11),
TO_SIGNED(-26,11),
TO_SIGNED(21,11),
TO_SIGNED(68,11),
TO_SIGNED(115,11),
TO_SIGNED(161,11),
TO_SIGNED(207,11),
TO_SIGNED(251,11),
TO_SIGNED(295,11),
TO_SIGNED(338,11),
TO_SIGNED(379,11),
TO_SIGNED(419,11),
TO_SIGNED(457,11),
TO_SIGNED(493,11),
TO_SIGNED(528,11),
TO_SIGNED(560,11),
TO_SIGNED(590,11),
TO_SIGNED(618,11),
TO_SIGNED(644,11),
TO_SIGNED(666,11),
TO_SIGNED(687,11),
TO_SIGNED(704,11),
TO_SIGNED(719,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(671,11),
TO_SIGNED(648,11),
TO_SIGNED(624,11),
TO_SIGNED(596,11),
TO_SIGNED(567,11),
TO_SIGNED(535,11),
TO_SIGNED(501,11),
TO_SIGNED(465,11),
TO_SIGNED(427,11),
TO_SIGNED(387,11),
TO_SIGNED(346,11),
TO_SIGNED(304,11),
TO_SIGNED(261,11),
TO_SIGNED(216,11),
TO_SIGNED(171,11),
TO_SIGNED(124,11),
TO_SIGNED(78,11),
TO_SIGNED(31,11),
TO_SIGNED(-16,11),
TO_SIGNED(-63,11),
TO_SIGNED(-110,11),
TO_SIGNED(-156,11),
TO_SIGNED(-202,11),
TO_SIGNED(-246,11),
TO_SIGNED(-290,11),
TO_SIGNED(-333,11),
TO_SIGNED(-375,11),
TO_SIGNED(-415,11),
TO_SIGNED(-453,11),
TO_SIGNED(-489,11),
TO_SIGNED(-524,11),
TO_SIGNED(-557,11),
TO_SIGNED(-587,11),
TO_SIGNED(-615,11),
TO_SIGNED(-641,11),
TO_SIGNED(-664,11),
TO_SIGNED(-685,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-730,11),
TO_SIGNED(-739,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-693,11),
TO_SIGNED(-673,11),
TO_SIGNED(-651,11),
TO_SIGNED(-627,11),
TO_SIGNED(-599,11),
TO_SIGNED(-570,11),
TO_SIGNED(-538,11),
TO_SIGNED(-505,11),
TO_SIGNED(-469,11),
TO_SIGNED(-431,11),
TO_SIGNED(-392,11),
TO_SIGNED(-351,11),
TO_SIGNED(-309,11),
TO_SIGNED(-266,11),
TO_SIGNED(-221,11),
TO_SIGNED(-176,11),
TO_SIGNED(-130,11),
TO_SIGNED(-83,11),
TO_SIGNED(-36,11),
TO_SIGNED(11,11),
TO_SIGNED(58,11),
TO_SIGNED(104,11),
TO_SIGNED(151,11),
TO_SIGNED(196,11),
TO_SIGNED(241,11),
TO_SIGNED(285,11),
TO_SIGNED(328,11),
TO_SIGNED(370,11),
TO_SIGNED(410,11),
TO_SIGNED(449,11),
TO_SIGNED(485,11),
TO_SIGNED(520,11),
TO_SIGNED(553,11),
TO_SIGNED(584,11),
TO_SIGNED(612,11),
TO_SIGNED(638,11),
TO_SIGNED(661,11),
TO_SIGNED(682,11),
TO_SIGNED(700,11),
TO_SIGNED(716,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(725,11),
TO_SIGNED(711,11),
TO_SIGNED(695,11),
TO_SIGNED(675,11),
TO_SIGNED(654,11),
TO_SIGNED(629,11),
TO_SIGNED(603,11),
TO_SIGNED(574,11),
TO_SIGNED(542,11),
TO_SIGNED(509,11),
TO_SIGNED(473,11),
TO_SIGNED(436,11),
TO_SIGNED(397,11),
TO_SIGNED(356,11),
TO_SIGNED(314,11),
TO_SIGNED(271,11),
TO_SIGNED(226,11),
TO_SIGNED(181,11),
TO_SIGNED(135,11),
TO_SIGNED(88,11),
TO_SIGNED(42,11),
TO_SIGNED(-5,11),
TO_SIGNED(-52,11),
TO_SIGNED(-99,11),
TO_SIGNED(-145,11),
TO_SIGNED(-191,11),
TO_SIGNED(-236,11),
TO_SIGNED(-280,11),
TO_SIGNED(-323,11),
TO_SIGNED(-365,11),
TO_SIGNED(-406,11),
TO_SIGNED(-444,11),
TO_SIGNED(-481,11),
TO_SIGNED(-516,11),
TO_SIGNED(-549,11),
TO_SIGNED(-580,11),
TO_SIGNED(-609,11),
TO_SIGNED(-635,11),
TO_SIGNED(-659,11),
TO_SIGNED(-680,11),
TO_SIGNED(-699,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-736,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-678,11),
TO_SIGNED(-656,11),
TO_SIGNED(-632,11),
TO_SIGNED(-606,11),
TO_SIGNED(-577,11),
TO_SIGNED(-546,11),
TO_SIGNED(-512,11),
TO_SIGNED(-477,11),
TO_SIGNED(-440,11),
TO_SIGNED(-401,11),
TO_SIGNED(-361,11),
TO_SIGNED(-319,11),
TO_SIGNED(-275,11),
TO_SIGNED(-231,11),
TO_SIGNED(-186,11),
TO_SIGNED(-140,11),
TO_SIGNED(-94,11),
TO_SIGNED(-47,11),
TO_SIGNED(0,11),
TO_SIGNED(47,11),
TO_SIGNED(94,11),
TO_SIGNED(140,11),
TO_SIGNED(186,11),
TO_SIGNED(231,11),
TO_SIGNED(275,11),
TO_SIGNED(319,11),
TO_SIGNED(361,11),
TO_SIGNED(401,11),
TO_SIGNED(440,11),
TO_SIGNED(477,11),
TO_SIGNED(512,11),
TO_SIGNED(546,11),
TO_SIGNED(577,11),
TO_SIGNED(606,11),
TO_SIGNED(632,11),
TO_SIGNED(656,11),
TO_SIGNED(678,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(736,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(699,11),
TO_SIGNED(680,11),
TO_SIGNED(659,11),
TO_SIGNED(635,11),
TO_SIGNED(609,11),
TO_SIGNED(580,11),
TO_SIGNED(549,11),
TO_SIGNED(516,11),
TO_SIGNED(481,11),
TO_SIGNED(444,11),
TO_SIGNED(406,11),
TO_SIGNED(365,11),
TO_SIGNED(323,11),
TO_SIGNED(280,11),
TO_SIGNED(236,11),
TO_SIGNED(191,11),
TO_SIGNED(145,11),
TO_SIGNED(99,11),
TO_SIGNED(52,11),
TO_SIGNED(5,11),
TO_SIGNED(-42,11),
TO_SIGNED(-88,11),
TO_SIGNED(-135,11),
TO_SIGNED(-181,11),
TO_SIGNED(-226,11),
TO_SIGNED(-271,11),
TO_SIGNED(-314,11),
TO_SIGNED(-356,11),
TO_SIGNED(-397,11),
TO_SIGNED(-436,11),
TO_SIGNED(-473,11),
TO_SIGNED(-509,11),
TO_SIGNED(-542,11),
TO_SIGNED(-574,11),
TO_SIGNED(-603,11),
TO_SIGNED(-629,11),
TO_SIGNED(-654,11),
TO_SIGNED(-675,11),
TO_SIGNED(-695,11),
TO_SIGNED(-711,11),
TO_SIGNED(-725,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-716,11),
TO_SIGNED(-700,11),
TO_SIGNED(-682,11),
TO_SIGNED(-661,11),
TO_SIGNED(-638,11),
TO_SIGNED(-612,11),
TO_SIGNED(-584,11),
TO_SIGNED(-553,11),
TO_SIGNED(-520,11),
TO_SIGNED(-485,11),
TO_SIGNED(-449,11),
TO_SIGNED(-410,11),
TO_SIGNED(-370,11),
TO_SIGNED(-328,11),
TO_SIGNED(-285,11),
TO_SIGNED(-241,11),
TO_SIGNED(-196,11),
TO_SIGNED(-151,11),
TO_SIGNED(-104,11),
TO_SIGNED(-58,11),
TO_SIGNED(-11,11),
TO_SIGNED(36,11),
TO_SIGNED(83,11),
TO_SIGNED(130,11),
TO_SIGNED(176,11),
TO_SIGNED(221,11),
TO_SIGNED(266,11),
TO_SIGNED(309,11),
TO_SIGNED(351,11),
TO_SIGNED(392,11),
TO_SIGNED(431,11),
TO_SIGNED(469,11),
TO_SIGNED(505,11),
TO_SIGNED(538,11),
TO_SIGNED(570,11),
TO_SIGNED(599,11),
TO_SIGNED(627,11),
TO_SIGNED(651,11),
TO_SIGNED(673,11),
TO_SIGNED(693,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(739,11),
TO_SIGNED(730,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(685,11),
TO_SIGNED(664,11),
TO_SIGNED(641,11),
TO_SIGNED(615,11),
TO_SIGNED(587,11),
TO_SIGNED(557,11),
TO_SIGNED(524,11),
TO_SIGNED(489,11),
TO_SIGNED(453,11),
TO_SIGNED(415,11),
TO_SIGNED(375,11),
TO_SIGNED(333,11),
TO_SIGNED(290,11),
TO_SIGNED(246,11),
TO_SIGNED(202,11),
TO_SIGNED(156,11),
TO_SIGNED(110,11),
TO_SIGNED(63,11),
TO_SIGNED(16,11),
TO_SIGNED(-31,11),
TO_SIGNED(-78,11),
TO_SIGNED(-124,11),
TO_SIGNED(-171,11),
TO_SIGNED(-216,11),
TO_SIGNED(-261,11),
TO_SIGNED(-304,11),
TO_SIGNED(-346,11),
TO_SIGNED(-387,11),
TO_SIGNED(-427,11),
TO_SIGNED(-465,11),
TO_SIGNED(-501,11),
TO_SIGNED(-535,11),
TO_SIGNED(-567,11),
TO_SIGNED(-596,11),
TO_SIGNED(-624,11),
TO_SIGNED(-648,11),
TO_SIGNED(-671,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-719,11),
TO_SIGNED(-704,11),
TO_SIGNED(-687,11),
TO_SIGNED(-666,11),
TO_SIGNED(-644,11),
TO_SIGNED(-618,11),
TO_SIGNED(-590,11),
TO_SIGNED(-560,11),
TO_SIGNED(-528,11),
TO_SIGNED(-493,11),
TO_SIGNED(-457,11),
TO_SIGNED(-419,11),
TO_SIGNED(-379,11),
TO_SIGNED(-338,11),
TO_SIGNED(-295,11),
TO_SIGNED(-251,11),
TO_SIGNED(-207,11),
TO_SIGNED(-161,11),
TO_SIGNED(-115,11),
TO_SIGNED(-68,11),
TO_SIGNED(-21,11),
TO_SIGNED(26,11),
TO_SIGNED(73,11),
TO_SIGNED(119,11),
TO_SIGNED(165,11),
TO_SIGNED(211,11),
TO_SIGNED(256,11),
TO_SIGNED(299,11),
TO_SIGNED(342,11),
TO_SIGNED(383,11),
TO_SIGNED(422,11),
TO_SIGNED(460,11),
TO_SIGNED(497,11),
TO_SIGNED(531,11),
TO_SIGNED(563,11),
TO_SIGNED(593,11),
TO_SIGNED(621,11),
TO_SIGNED(646,11),
TO_SIGNED(668,11),
TO_SIGNED(688,11),
TO_SIGNED(706,11),
TO_SIGNED(720,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(721,11),
TO_SIGNED(706,11),
TO_SIGNED(689,11),
TO_SIGNED(669,11),
TO_SIGNED(646,11),
TO_SIGNED(621,11),
TO_SIGNED(594,11),
TO_SIGNED(564,11),
TO_SIGNED(532,11),
TO_SIGNED(497,11),
TO_SIGNED(461,11),
TO_SIGNED(423,11),
TO_SIGNED(384,11),
TO_SIGNED(343,11),
TO_SIGNED(300,11),
TO_SIGNED(257,11),
TO_SIGNED(212,11),
TO_SIGNED(166,11),
TO_SIGNED(120,11),
TO_SIGNED(74,11),
TO_SIGNED(27,11),
TO_SIGNED(-20,11),
TO_SIGNED(-67,11),
TO_SIGNED(-114,11),
TO_SIGNED(-160,11),
TO_SIGNED(-206,11),
TO_SIGNED(-250,11),
TO_SIGNED(-294,11),
TO_SIGNED(-337,11),
TO_SIGNED(-378,11),
TO_SIGNED(-418,11),
TO_SIGNED(-456,11),
TO_SIGNED(-493,11),
TO_SIGNED(-527,11),
TO_SIGNED(-559,11),
TO_SIGNED(-590,11),
TO_SIGNED(-618,11),
TO_SIGNED(-643,11),
TO_SIGNED(-666,11),
TO_SIGNED(-686,11),
TO_SIGNED(-704,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-733,11),
TO_SIGNED(-722,11),
TO_SIGNED(-708,11),
TO_SIGNED(-691,11),
TO_SIGNED(-671,11),
TO_SIGNED(-649,11),
TO_SIGNED(-624,11),
TO_SIGNED(-597,11),
TO_SIGNED(-567,11),
TO_SIGNED(-535,11),
TO_SIGNED(-501,11),
TO_SIGNED(-466,11),
TO_SIGNED(-428,11),
TO_SIGNED(-388,11),
TO_SIGNED(-347,11),
TO_SIGNED(-305,11),
TO_SIGNED(-262,11),
TO_SIGNED(-217,11),
TO_SIGNED(-172,11),
TO_SIGNED(-125,11),
TO_SIGNED(-79,11),
TO_SIGNED(-32,11),
TO_SIGNED(15,11),
TO_SIGNED(62,11),
TO_SIGNED(109,11),
TO_SIGNED(155,11),
TO_SIGNED(201,11),
TO_SIGNED(245,11),
TO_SIGNED(289,11),
TO_SIGNED(332,11),
TO_SIGNED(374,11),
TO_SIGNED(414,11),
TO_SIGNED(452,11),
TO_SIGNED(489,11),
TO_SIGNED(523,11),
TO_SIGNED(556,11),
TO_SIGNED(586,11),
TO_SIGNED(615,11),
TO_SIGNED(640,11),
TO_SIGNED(663,11),
TO_SIGNED(684,11),
TO_SIGNED(702,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(710,11),
TO_SIGNED(693,11),
TO_SIGNED(674,11),
TO_SIGNED(652,11),
TO_SIGNED(627,11),
TO_SIGNED(600,11),
TO_SIGNED(571,11),
TO_SIGNED(539,11),
TO_SIGNED(505,11),
TO_SIGNED(470,11),
TO_SIGNED(432,11),
TO_SIGNED(393,11),
TO_SIGNED(352,11),
TO_SIGNED(310,11),
TO_SIGNED(267,11),
TO_SIGNED(222,11),
TO_SIGNED(177,11),
TO_SIGNED(131,11),
TO_SIGNED(84,11),
TO_SIGNED(37,11),
TO_SIGNED(-10,11),
TO_SIGNED(-57,11),
TO_SIGNED(-103,11),
TO_SIGNED(-150,11),
TO_SIGNED(-195,11),
TO_SIGNED(-240,11),
TO_SIGNED(-284,11),
TO_SIGNED(-327,11),
TO_SIGNED(-369,11),
TO_SIGNED(-409,11),
TO_SIGNED(-448,11),
TO_SIGNED(-485,11),
TO_SIGNED(-519,11),
TO_SIGNED(-552,11),
TO_SIGNED(-583,11),
TO_SIGNED(-611,11),
TO_SIGNED(-637,11),
TO_SIGNED(-661,11),
TO_SIGNED(-682,11),
TO_SIGNED(-700,11),
TO_SIGNED(-716,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-725,11),
TO_SIGNED(-711,11),
TO_SIGNED(-695,11),
TO_SIGNED(-676,11),
TO_SIGNED(-654,11),
TO_SIGNED(-630,11),
TO_SIGNED(-603,11),
TO_SIGNED(-574,11),
TO_SIGNED(-543,11),
TO_SIGNED(-509,11),
TO_SIGNED(-474,11),
TO_SIGNED(-437,11),
TO_SIGNED(-397,11),
TO_SIGNED(-357,11),
TO_SIGNED(-315,11),
TO_SIGNED(-272,11),
TO_SIGNED(-227,11),
TO_SIGNED(-182,11),
TO_SIGNED(-136,11),
TO_SIGNED(-90,11),
TO_SIGNED(-43,11),
TO_SIGNED(4,11),
TO_SIGNED(51,11),
TO_SIGNED(98,11),
TO_SIGNED(144,11),
TO_SIGNED(190,11),
TO_SIGNED(235,11),
TO_SIGNED(279,11),
TO_SIGNED(323,11),
TO_SIGNED(364,11),
TO_SIGNED(405,11),
TO_SIGNED(443,11),
TO_SIGNED(480,11),
TO_SIGNED(516,11),
TO_SIGNED(549,11),
TO_SIGNED(580,11),
TO_SIGNED(608,11),
TO_SIGNED(635,11),
TO_SIGNED(658,11),
TO_SIGNED(680,11),
TO_SIGNED(698,11),
TO_SIGNED(714,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(713,11),
TO_SIGNED(697,11),
TO_SIGNED(678,11),
TO_SIGNED(657,11),
TO_SIGNED(633,11),
TO_SIGNED(606,11),
TO_SIGNED(578,11),
TO_SIGNED(547,11),
TO_SIGNED(513,11),
TO_SIGNED(478,11),
TO_SIGNED(441,11),
TO_SIGNED(402,11),
TO_SIGNED(362,11),
TO_SIGNED(320,11),
TO_SIGNED(276,11),
TO_SIGNED(232,11),
TO_SIGNED(187,11),
TO_SIGNED(141,11),
TO_SIGNED(95,11),
TO_SIGNED(48,11),
TO_SIGNED(1,11),
TO_SIGNED(-46,11),
TO_SIGNED(-93,11),
TO_SIGNED(-139,11),
TO_SIGNED(-185,11),
TO_SIGNED(-230,11),
TO_SIGNED(-275,11),
TO_SIGNED(-318,11),
TO_SIGNED(-360,11),
TO_SIGNED(-400,11),
TO_SIGNED(-439,11),
TO_SIGNED(-476,11),
TO_SIGNED(-512,11),
TO_SIGNED(-545,11),
TO_SIGNED(-576,11),
TO_SIGNED(-605,11),
TO_SIGNED(-632,11),
TO_SIGNED(-656,11),
TO_SIGNED(-677,11),
TO_SIGNED(-696,11),
TO_SIGNED(-712,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-715,11),
TO_SIGNED(-699,11),
TO_SIGNED(-681,11),
TO_SIGNED(-659,11),
TO_SIGNED(-636,11),
TO_SIGNED(-610,11),
TO_SIGNED(-581,11),
TO_SIGNED(-550,11),
TO_SIGNED(-517,11),
TO_SIGNED(-482,11),
TO_SIGNED(-445,11),
TO_SIGNED(-406,11),
TO_SIGNED(-366,11),
TO_SIGNED(-324,11),
TO_SIGNED(-281,11),
TO_SIGNED(-237,11),
TO_SIGNED(-192,11),
TO_SIGNED(-147,11),
TO_SIGNED(-100,11),
TO_SIGNED(-53,11),
TO_SIGNED(-6,11),
TO_SIGNED(41,11),
TO_SIGNED(87,11),
TO_SIGNED(134,11),
TO_SIGNED(180,11),
TO_SIGNED(225,11),
TO_SIGNED(270,11),
TO_SIGNED(313,11),
TO_SIGNED(355,11),
TO_SIGNED(396,11),
TO_SIGNED(435,11),
TO_SIGNED(472,11),
TO_SIGNED(508,11),
TO_SIGNED(541,11),
TO_SIGNED(573,11),
TO_SIGNED(602,11),
TO_SIGNED(629,11),
TO_SIGNED(653,11),
TO_SIGNED(675,11),
TO_SIGNED(694,11),
TO_SIGNED(711,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(729,11),
TO_SIGNED(716,11),
TO_SIGNED(701,11),
TO_SIGNED(683,11),
TO_SIGNED(662,11),
TO_SIGNED(639,11),
TO_SIGNED(613,11),
TO_SIGNED(584,11),
TO_SIGNED(554,11),
TO_SIGNED(521,11),
TO_SIGNED(486,11),
TO_SIGNED(449,11),
TO_SIGNED(411,11),
TO_SIGNED(371,11),
TO_SIGNED(329,11),
TO_SIGNED(286,11),
TO_SIGNED(242,11),
TO_SIGNED(197,11),
TO_SIGNED(152,11),
TO_SIGNED(105,11),
TO_SIGNED(59,11),
TO_SIGNED(12,11),
TO_SIGNED(-35,11),
TO_SIGNED(-82,11),
TO_SIGNED(-129,11),
TO_SIGNED(-175,11),
TO_SIGNED(-220,11),
TO_SIGNED(-265,11),
TO_SIGNED(-308,11),
TO_SIGNED(-350,11),
TO_SIGNED(-391,11),
TO_SIGNED(-430,11),
TO_SIGNED(-468,11),
TO_SIGNED(-504,11),
TO_SIGNED(-538,11),
TO_SIGNED(-569,11),
TO_SIGNED(-599,11),
TO_SIGNED(-626,11),
TO_SIGNED(-651,11),
TO_SIGNED(-673,11),
TO_SIGNED(-692,11),
TO_SIGNED(-709,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-685,11),
TO_SIGNED(-664,11),
TO_SIGNED(-641,11),
TO_SIGNED(-616,11),
TO_SIGNED(-588,11),
TO_SIGNED(-557,11),
TO_SIGNED(-525,11),
TO_SIGNED(-490,11),
TO_SIGNED(-454,11),
TO_SIGNED(-415,11),
TO_SIGNED(-375,11),
TO_SIGNED(-334,11),
TO_SIGNED(-291,11),
TO_SIGNED(-247,11),
TO_SIGNED(-203,11),
TO_SIGNED(-157,11),
TO_SIGNED(-111,11),
TO_SIGNED(-64,11),
TO_SIGNED(-17,11),
TO_SIGNED(30,11),
TO_SIGNED(77,11),
TO_SIGNED(123,11),
TO_SIGNED(169,11),
TO_SIGNED(215,11),
TO_SIGNED(260,11),
TO_SIGNED(303,11),
TO_SIGNED(345,11),
TO_SIGNED(387,11),
TO_SIGNED(426,11),
TO_SIGNED(464,11),
TO_SIGNED(500,11),
TO_SIGNED(534,11),
TO_SIGNED(566,11),
TO_SIGNED(596,11),
TO_SIGNED(623,11),
TO_SIGNED(648,11),
TO_SIGNED(670,11),
TO_SIGNED(690,11),
TO_SIGNED(707,11),
TO_SIGNED(721,11),
TO_SIGNED(733,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(705,11),
TO_SIGNED(687,11),
TO_SIGNED(667,11),
TO_SIGNED(644,11),
TO_SIGNED(619,11),
TO_SIGNED(591,11),
TO_SIGNED(561,11),
TO_SIGNED(529,11),
TO_SIGNED(494,11),
TO_SIGNED(458,11),
TO_SIGNED(420,11),
TO_SIGNED(380,11),
TO_SIGNED(339,11),
TO_SIGNED(296,11),
TO_SIGNED(252,11),
TO_SIGNED(208,11),
TO_SIGNED(162,11),
TO_SIGNED(116,11),
TO_SIGNED(69,11),
TO_SIGNED(22,11),
TO_SIGNED(-25,11),
TO_SIGNED(-71,11),
TO_SIGNED(-118,11),
TO_SIGNED(-164,11),
TO_SIGNED(-210,11),
TO_SIGNED(-255,11),
TO_SIGNED(-298,11),
TO_SIGNED(-341,11),
TO_SIGNED(-382,11),
TO_SIGNED(-422,11),
TO_SIGNED(-460,11),
TO_SIGNED(-496,11),
TO_SIGNED(-530,11),
TO_SIGNED(-562,11),
TO_SIGNED(-592,11),
TO_SIGNED(-620,11),
TO_SIGNED(-645,11),
TO_SIGNED(-668,11),
TO_SIGNED(-688,11),
TO_SIGNED(-705,11),
TO_SIGNED(-720,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-721,11),
TO_SIGNED(-706,11),
TO_SIGNED(-689,11),
TO_SIGNED(-669,11),
TO_SIGNED(-647,11),
TO_SIGNED(-622,11),
TO_SIGNED(-594,11),
TO_SIGNED(-564,11),
TO_SIGNED(-532,11),
TO_SIGNED(-498,11),
TO_SIGNED(-462,11),
TO_SIGNED(-424,11),
TO_SIGNED(-385,11),
TO_SIGNED(-344,11),
TO_SIGNED(-301,11),
TO_SIGNED(-258,11),
TO_SIGNED(-213,11),
TO_SIGNED(-167,11),
TO_SIGNED(-121,11),
TO_SIGNED(-75,11),
TO_SIGNED(-28,11),
TO_SIGNED(19,11),
TO_SIGNED(66,11),
TO_SIGNED(113,11),
TO_SIGNED(159,11),
TO_SIGNED(205,11),
TO_SIGNED(249,11),
TO_SIGNED(293,11),
TO_SIGNED(336,11),
TO_SIGNED(377,11),
TO_SIGNED(417,11),
TO_SIGNED(455,11),
TO_SIGNED(492,11),
TO_SIGNED(526,11),
TO_SIGNED(559,11),
TO_SIGNED(589,11),
TO_SIGNED(617,11),
TO_SIGNED(642,11),
TO_SIGNED(665,11),
TO_SIGNED(686,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(708,11),
TO_SIGNED(691,11),
TO_SIGNED(672,11),
TO_SIGNED(650,11),
TO_SIGNED(625,11),
TO_SIGNED(598,11),
TO_SIGNED(568,11),
TO_SIGNED(536,11),
TO_SIGNED(502,11),
TO_SIGNED(466,11),
TO_SIGNED(429,11),
TO_SIGNED(389,11),
TO_SIGNED(348,11),
TO_SIGNED(306,11),
TO_SIGNED(263,11),
TO_SIGNED(218,11),
TO_SIGNED(173,11),
TO_SIGNED(127,11),
TO_SIGNED(80,11),
TO_SIGNED(33,11),
TO_SIGNED(-14,11),
TO_SIGNED(-61,11),
TO_SIGNED(-108,11),
TO_SIGNED(-154,11),
TO_SIGNED(-200,11),
TO_SIGNED(-244,11),
TO_SIGNED(-288,11),
TO_SIGNED(-331,11),
TO_SIGNED(-373,11),
TO_SIGNED(-413,11),
TO_SIGNED(-451,11),
TO_SIGNED(-488,11),
TO_SIGNED(-523,11),
TO_SIGNED(-555,11),
TO_SIGNED(-586,11),
TO_SIGNED(-614,11),
TO_SIGNED(-640,11),
TO_SIGNED(-663,11),
TO_SIGNED(-684,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-729,11),
TO_SIGNED(-739,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-710,11),
TO_SIGNED(-693,11),
TO_SIGNED(-674,11),
TO_SIGNED(-652,11),
TO_SIGNED(-628,11),
TO_SIGNED(-601,11),
TO_SIGNED(-571,11),
TO_SIGNED(-540,11),
TO_SIGNED(-506,11),
TO_SIGNED(-471,11),
TO_SIGNED(-433,11),
TO_SIGNED(-394,11),
TO_SIGNED(-353,11),
TO_SIGNED(-311,11),
TO_SIGNED(-268,11),
TO_SIGNED(-223,11),
TO_SIGNED(-178,11),
TO_SIGNED(-132,11),
TO_SIGNED(-85,11),
TO_SIGNED(-38,11),
TO_SIGNED(9,11),
TO_SIGNED(56,11),
TO_SIGNED(102,11),
TO_SIGNED(149,11),
TO_SIGNED(194,11),
TO_SIGNED(239,11),
TO_SIGNED(283,11),
TO_SIGNED(326,11),
TO_SIGNED(368,11),
TO_SIGNED(408,11),
TO_SIGNED(447,11),
TO_SIGNED(484,11),
TO_SIGNED(519,11),
TO_SIGNED(552,11),
TO_SIGNED(582,11),
TO_SIGNED(611,11),
TO_SIGNED(637,11),
TO_SIGNED(660,11),
TO_SIGNED(681,11),
TO_SIGNED(700,11),
TO_SIGNED(715,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(736,11),
TO_SIGNED(725,11),
TO_SIGNED(712,11),
TO_SIGNED(695,11),
TO_SIGNED(676,11),
TO_SIGNED(655,11),
TO_SIGNED(631,11),
TO_SIGNED(604,11),
TO_SIGNED(575,11),
TO_SIGNED(544,11),
TO_SIGNED(510,11),
TO_SIGNED(475,11),
TO_SIGNED(437,11),
TO_SIGNED(398,11),
TO_SIGNED(358,11),
TO_SIGNED(316,11),
TO_SIGNED(273,11),
TO_SIGNED(228,11),
TO_SIGNED(183,11),
TO_SIGNED(137,11),
TO_SIGNED(91,11),
TO_SIGNED(44,11),
TO_SIGNED(-3,11),
TO_SIGNED(-50,11),
TO_SIGNED(-97,11),
TO_SIGNED(-143,11),
TO_SIGNED(-189,11),
TO_SIGNED(-234,11),
TO_SIGNED(-278,11),
TO_SIGNED(-322,11),
TO_SIGNED(-363,11),
TO_SIGNED(-404,11),
TO_SIGNED(-443,11),
TO_SIGNED(-480,11),
TO_SIGNED(-515,11),
TO_SIGNED(-548,11),
TO_SIGNED(-579,11),
TO_SIGNED(-608,11),
TO_SIGNED(-634,11),
TO_SIGNED(-658,11),
TO_SIGNED(-679,11),
TO_SIGNED(-698,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-679,11),
TO_SIGNED(-657,11),
TO_SIGNED(-633,11),
TO_SIGNED(-607,11),
TO_SIGNED(-578,11),
TO_SIGNED(-547,11),
TO_SIGNED(-514,11),
TO_SIGNED(-479,11),
TO_SIGNED(-442,11),
TO_SIGNED(-403,11),
TO_SIGNED(-362,11),
TO_SIGNED(-321,11),
TO_SIGNED(-277,11),
TO_SIGNED(-233,11),
TO_SIGNED(-188,11),
TO_SIGNED(-142,11),
TO_SIGNED(-96,11),
TO_SIGNED(-49,11),
TO_SIGNED(-2,11),
TO_SIGNED(45,11),
TO_SIGNED(92,11),
TO_SIGNED(138,11),
TO_SIGNED(184,11),
TO_SIGNED(229,11),
TO_SIGNED(274,11),
TO_SIGNED(317,11),
TO_SIGNED(359,11),
TO_SIGNED(399,11),
TO_SIGNED(438,11),
TO_SIGNED(476,11),
TO_SIGNED(511,11),
TO_SIGNED(544,11),
TO_SIGNED(576,11),
TO_SIGNED(605,11),
TO_SIGNED(631,11),
TO_SIGNED(655,11),
TO_SIGNED(677,11),
TO_SIGNED(696,11),
TO_SIGNED(712,11),
TO_SIGNED(725,11),
TO_SIGNED(736,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(715,11),
TO_SIGNED(699,11),
TO_SIGNED(681,11),
TO_SIGNED(660,11),
TO_SIGNED(636,11),
TO_SIGNED(610,11),
TO_SIGNED(582,11),
TO_SIGNED(551,11),
TO_SIGNED(518,11),
TO_SIGNED(483,11),
TO_SIGNED(446,11),
TO_SIGNED(407,11),
TO_SIGNED(367,11),
TO_SIGNED(325,11),
TO_SIGNED(282,11),
TO_SIGNED(238,11),
TO_SIGNED(193,11),
TO_SIGNED(148,11),
TO_SIGNED(101,11),
TO_SIGNED(54,11),
TO_SIGNED(7,11),
TO_SIGNED(-40,11),
TO_SIGNED(-86,11),
TO_SIGNED(-133,11),
TO_SIGNED(-179,11),
TO_SIGNED(-224,11),
TO_SIGNED(-269,11),
TO_SIGNED(-312,11),
TO_SIGNED(-354,11),
TO_SIGNED(-395,11),
TO_SIGNED(-434,11),
TO_SIGNED(-471,11),
TO_SIGNED(-507,11),
TO_SIGNED(-541,11),
TO_SIGNED(-572,11),
TO_SIGNED(-601,11),
TO_SIGNED(-628,11),
TO_SIGNED(-653,11),
TO_SIGNED(-675,11),
TO_SIGNED(-694,11),
TO_SIGNED(-710,11),
TO_SIGNED(-724,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-701,11),
TO_SIGNED(-683,11),
TO_SIGNED(-662,11),
TO_SIGNED(-639,11),
TO_SIGNED(-613,11),
TO_SIGNED(-585,11),
TO_SIGNED(-554,11),
TO_SIGNED(-522,11),
TO_SIGNED(-487,11),
TO_SIGNED(-450,11),
TO_SIGNED(-412,11),
TO_SIGNED(-372,11),
TO_SIGNED(-330,11),
TO_SIGNED(-287,11),
TO_SIGNED(-243,11),
TO_SIGNED(-198,11),
TO_SIGNED(-153,11),
TO_SIGNED(-106,11),
TO_SIGNED(-60,11),
TO_SIGNED(-13,11),
TO_SIGNED(34,11),
TO_SIGNED(81,11),
TO_SIGNED(128,11),
TO_SIGNED(174,11),
TO_SIGNED(219,11),
TO_SIGNED(264,11),
TO_SIGNED(307,11),
TO_SIGNED(349,11),
TO_SIGNED(390,11),
TO_SIGNED(430,11),
TO_SIGNED(467,11),
TO_SIGNED(503,11),
TO_SIGNED(537,11),
TO_SIGNED(569,11),
TO_SIGNED(598,11),
TO_SIGNED(625,11),
TO_SIGNED(650,11),
TO_SIGNED(672,11),
TO_SIGNED(692,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(730,11),
TO_SIGNED(718,11),
TO_SIGNED(703,11),
TO_SIGNED(685,11),
TO_SIGNED(665,11),
TO_SIGNED(642,11),
TO_SIGNED(616,11),
TO_SIGNED(588,11),
TO_SIGNED(558,11),
TO_SIGNED(526,11),
TO_SIGNED(491,11),
TO_SIGNED(455,11),
TO_SIGNED(416,11),
TO_SIGNED(376,11),
TO_SIGNED(335,11),
TO_SIGNED(292,11),
TO_SIGNED(248,11),
TO_SIGNED(204,11),
TO_SIGNED(158,11),
TO_SIGNED(112,11),
TO_SIGNED(65,11),
TO_SIGNED(18,11),
TO_SIGNED(-29,11),
TO_SIGNED(-76,11),
TO_SIGNED(-122,11),
TO_SIGNED(-168,11),
TO_SIGNED(-214,11),
TO_SIGNED(-259,11),
TO_SIGNED(-302,11),
TO_SIGNED(-345,11),
TO_SIGNED(-386,11),
TO_SIGNED(-425,11),
TO_SIGNED(-463,11),
TO_SIGNED(-499,11),
TO_SIGNED(-533,11),
TO_SIGNED(-565,11),
TO_SIGNED(-595,11),
TO_SIGNED(-622,11),
TO_SIGNED(-647,11),
TO_SIGNED(-670,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-721,11),
TO_SIGNED(-733,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-720,11),
TO_SIGNED(-705,11),
TO_SIGNED(-688,11),
TO_SIGNED(-667,11),
TO_SIGNED(-645,11),
TO_SIGNED(-619,11),
TO_SIGNED(-592,11),
TO_SIGNED(-562,11),
TO_SIGNED(-529,11),
TO_SIGNED(-495,11),
TO_SIGNED(-459,11),
TO_SIGNED(-421,11),
TO_SIGNED(-381,11),
TO_SIGNED(-340,11),
TO_SIGNED(-297,11),
TO_SIGNED(-254,11),
TO_SIGNED(-209,11),
TO_SIGNED(-163,11),
TO_SIGNED(-117,11),
TO_SIGNED(-70,11),
TO_SIGNED(-24,11),
TO_SIGNED(24,11),
TO_SIGNED(70,11),
TO_SIGNED(117,11),
TO_SIGNED(163,11),
TO_SIGNED(209,11),
TO_SIGNED(254,11),
TO_SIGNED(297,11),
TO_SIGNED(340,11),
TO_SIGNED(381,11),
TO_SIGNED(421,11),
TO_SIGNED(459,11),
TO_SIGNED(495,11),
TO_SIGNED(529,11),
TO_SIGNED(562,11),
TO_SIGNED(592,11),
TO_SIGNED(619,11),
TO_SIGNED(645,11),
TO_SIGNED(667,11),
TO_SIGNED(688,11),
TO_SIGNED(705,11),
TO_SIGNED(720,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(733,11),
TO_SIGNED(721,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(670,11),
TO_SIGNED(647,11),
TO_SIGNED(622,11),
TO_SIGNED(595,11),
TO_SIGNED(565,11),
TO_SIGNED(533,11),
TO_SIGNED(499,11),
TO_SIGNED(463,11),
TO_SIGNED(425,11),
TO_SIGNED(386,11),
TO_SIGNED(345,11),
TO_SIGNED(302,11),
TO_SIGNED(259,11),
TO_SIGNED(214,11),
TO_SIGNED(168,11),
TO_SIGNED(122,11),
TO_SIGNED(76,11),
TO_SIGNED(29,11),
TO_SIGNED(-18,11),
TO_SIGNED(-65,11),
TO_SIGNED(-112,11),
TO_SIGNED(-158,11),
TO_SIGNED(-204,11),
TO_SIGNED(-248,11),
TO_SIGNED(-292,11),
TO_SIGNED(-335,11),
TO_SIGNED(-376,11),
TO_SIGNED(-416,11),
TO_SIGNED(-455,11),
TO_SIGNED(-491,11),
TO_SIGNED(-526,11),
TO_SIGNED(-558,11),
TO_SIGNED(-588,11),
TO_SIGNED(-616,11),
TO_SIGNED(-642,11),
TO_SIGNED(-665,11),
TO_SIGNED(-685,11),
TO_SIGNED(-703,11),
TO_SIGNED(-718,11),
TO_SIGNED(-730,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-692,11),
TO_SIGNED(-672,11),
TO_SIGNED(-650,11),
TO_SIGNED(-625,11),
TO_SIGNED(-598,11),
TO_SIGNED(-569,11),
TO_SIGNED(-537,11),
TO_SIGNED(-503,11),
TO_SIGNED(-467,11),
TO_SIGNED(-430,11),
TO_SIGNED(-390,11),
TO_SIGNED(-349,11),
TO_SIGNED(-307,11),
TO_SIGNED(-264,11),
TO_SIGNED(-219,11),
TO_SIGNED(-174,11),
TO_SIGNED(-128,11),
TO_SIGNED(-81,11),
TO_SIGNED(-34,11),
TO_SIGNED(13,11),
TO_SIGNED(60,11),
TO_SIGNED(106,11),
TO_SIGNED(153,11),
TO_SIGNED(198,11),
TO_SIGNED(243,11),
TO_SIGNED(287,11),
TO_SIGNED(330,11),
TO_SIGNED(372,11),
TO_SIGNED(412,11),
TO_SIGNED(450,11),
TO_SIGNED(487,11),
TO_SIGNED(522,11),
TO_SIGNED(554,11),
TO_SIGNED(585,11),
TO_SIGNED(613,11),
TO_SIGNED(639,11),
TO_SIGNED(662,11),
TO_SIGNED(683,11),
TO_SIGNED(701,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(724,11),
TO_SIGNED(710,11),
TO_SIGNED(694,11),
TO_SIGNED(675,11),
TO_SIGNED(653,11),
TO_SIGNED(628,11),
TO_SIGNED(601,11),
TO_SIGNED(572,11),
TO_SIGNED(541,11),
TO_SIGNED(507,11),
TO_SIGNED(471,11),
TO_SIGNED(434,11),
TO_SIGNED(395,11),
TO_SIGNED(354,11),
TO_SIGNED(312,11),
TO_SIGNED(269,11),
TO_SIGNED(224,11),
TO_SIGNED(179,11),
TO_SIGNED(133,11),
TO_SIGNED(86,11),
TO_SIGNED(40,11),
TO_SIGNED(-7,11),
TO_SIGNED(-54,11),
TO_SIGNED(-101,11),
TO_SIGNED(-148,11),
TO_SIGNED(-193,11),
TO_SIGNED(-238,11),
TO_SIGNED(-282,11),
TO_SIGNED(-325,11),
TO_SIGNED(-367,11),
TO_SIGNED(-407,11),
TO_SIGNED(-446,11),
TO_SIGNED(-483,11),
TO_SIGNED(-518,11),
TO_SIGNED(-551,11),
TO_SIGNED(-582,11),
TO_SIGNED(-610,11),
TO_SIGNED(-636,11),
TO_SIGNED(-660,11),
TO_SIGNED(-681,11),
TO_SIGNED(-699,11),
TO_SIGNED(-715,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-736,11),
TO_SIGNED(-725,11),
TO_SIGNED(-712,11),
TO_SIGNED(-696,11),
TO_SIGNED(-677,11),
TO_SIGNED(-655,11),
TO_SIGNED(-631,11),
TO_SIGNED(-605,11),
TO_SIGNED(-576,11),
TO_SIGNED(-544,11),
TO_SIGNED(-511,11),
TO_SIGNED(-476,11),
TO_SIGNED(-438,11),
TO_SIGNED(-399,11),
TO_SIGNED(-359,11),
TO_SIGNED(-317,11),
TO_SIGNED(-274,11),
TO_SIGNED(-229,11),
TO_SIGNED(-184,11),
TO_SIGNED(-138,11),
TO_SIGNED(-92,11),
TO_SIGNED(-45,11),
TO_SIGNED(2,11),
TO_SIGNED(49,11),
TO_SIGNED(96,11),
TO_SIGNED(142,11),
TO_SIGNED(188,11),
TO_SIGNED(233,11),
TO_SIGNED(277,11),
TO_SIGNED(321,11),
TO_SIGNED(362,11),
TO_SIGNED(403,11),
TO_SIGNED(442,11),
TO_SIGNED(479,11),
TO_SIGNED(514,11),
TO_SIGNED(547,11),
TO_SIGNED(578,11),
TO_SIGNED(607,11),
TO_SIGNED(633,11),
TO_SIGNED(657,11),
TO_SIGNED(679,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(698,11),
TO_SIGNED(679,11),
TO_SIGNED(658,11),
TO_SIGNED(634,11),
TO_SIGNED(608,11),
TO_SIGNED(579,11),
TO_SIGNED(548,11),
TO_SIGNED(515,11),
TO_SIGNED(480,11),
TO_SIGNED(443,11),
TO_SIGNED(404,11),
TO_SIGNED(363,11),
TO_SIGNED(322,11),
TO_SIGNED(278,11),
TO_SIGNED(234,11),
TO_SIGNED(189,11),
TO_SIGNED(143,11),
TO_SIGNED(97,11),
TO_SIGNED(50,11),
TO_SIGNED(3,11),
TO_SIGNED(-44,11),
TO_SIGNED(-91,11),
TO_SIGNED(-137,11),
TO_SIGNED(-183,11),
TO_SIGNED(-228,11),
TO_SIGNED(-273,11),
TO_SIGNED(-316,11),
TO_SIGNED(-358,11),
TO_SIGNED(-398,11),
TO_SIGNED(-437,11),
TO_SIGNED(-475,11),
TO_SIGNED(-510,11),
TO_SIGNED(-544,11),
TO_SIGNED(-575,11),
TO_SIGNED(-604,11),
TO_SIGNED(-631,11),
TO_SIGNED(-655,11),
TO_SIGNED(-676,11),
TO_SIGNED(-695,11),
TO_SIGNED(-712,11),
TO_SIGNED(-725,11),
TO_SIGNED(-736,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-715,11),
TO_SIGNED(-700,11),
TO_SIGNED(-681,11),
TO_SIGNED(-660,11),
TO_SIGNED(-637,11),
TO_SIGNED(-611,11),
TO_SIGNED(-582,11),
TO_SIGNED(-552,11),
TO_SIGNED(-519,11),
TO_SIGNED(-484,11),
TO_SIGNED(-447,11),
TO_SIGNED(-408,11),
TO_SIGNED(-368,11),
TO_SIGNED(-326,11),
TO_SIGNED(-283,11),
TO_SIGNED(-239,11),
TO_SIGNED(-194,11),
TO_SIGNED(-149,11),
TO_SIGNED(-102,11),
TO_SIGNED(-56,11),
TO_SIGNED(-9,11),
TO_SIGNED(38,11),
TO_SIGNED(85,11),
TO_SIGNED(132,11),
TO_SIGNED(178,11),
TO_SIGNED(223,11),
TO_SIGNED(268,11),
TO_SIGNED(311,11),
TO_SIGNED(353,11),
TO_SIGNED(394,11),
TO_SIGNED(433,11),
TO_SIGNED(471,11),
TO_SIGNED(506,11),
TO_SIGNED(540,11),
TO_SIGNED(571,11),
TO_SIGNED(601,11),
TO_SIGNED(628,11),
TO_SIGNED(652,11),
TO_SIGNED(674,11),
TO_SIGNED(693,11),
TO_SIGNED(710,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(739,11),
TO_SIGNED(729,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(684,11),
TO_SIGNED(663,11),
TO_SIGNED(640,11),
TO_SIGNED(614,11),
TO_SIGNED(586,11),
TO_SIGNED(555,11),
TO_SIGNED(523,11),
TO_SIGNED(488,11),
TO_SIGNED(451,11),
TO_SIGNED(413,11),
TO_SIGNED(373,11),
TO_SIGNED(331,11),
TO_SIGNED(288,11),
TO_SIGNED(244,11),
TO_SIGNED(200,11),
TO_SIGNED(154,11),
TO_SIGNED(108,11),
TO_SIGNED(61,11),
TO_SIGNED(14,11),
TO_SIGNED(-33,11),
TO_SIGNED(-80,11),
TO_SIGNED(-127,11),
TO_SIGNED(-173,11),
TO_SIGNED(-218,11),
TO_SIGNED(-263,11),
TO_SIGNED(-306,11),
TO_SIGNED(-348,11),
TO_SIGNED(-389,11),
TO_SIGNED(-429,11),
TO_SIGNED(-466,11),
TO_SIGNED(-502,11),
TO_SIGNED(-536,11),
TO_SIGNED(-568,11),
TO_SIGNED(-598,11),
TO_SIGNED(-625,11),
TO_SIGNED(-650,11),
TO_SIGNED(-672,11),
TO_SIGNED(-691,11),
TO_SIGNED(-708,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-686,11),
TO_SIGNED(-665,11),
TO_SIGNED(-642,11),
TO_SIGNED(-617,11),
TO_SIGNED(-589,11),
TO_SIGNED(-559,11),
TO_SIGNED(-526,11),
TO_SIGNED(-492,11),
TO_SIGNED(-455,11),
TO_SIGNED(-417,11),
TO_SIGNED(-377,11),
TO_SIGNED(-336,11),
TO_SIGNED(-293,11),
TO_SIGNED(-249,11),
TO_SIGNED(-205,11),
TO_SIGNED(-159,11),
TO_SIGNED(-113,11),
TO_SIGNED(-66,11),
TO_SIGNED(-19,11),
TO_SIGNED(28,11),
TO_SIGNED(75,11),
TO_SIGNED(121,11),
TO_SIGNED(167,11),
TO_SIGNED(213,11),
TO_SIGNED(258,11),
TO_SIGNED(301,11),
TO_SIGNED(344,11),
TO_SIGNED(385,11),
TO_SIGNED(424,11),
TO_SIGNED(462,11),
TO_SIGNED(498,11),
TO_SIGNED(532,11),
TO_SIGNED(564,11),
TO_SIGNED(594,11),
TO_SIGNED(622,11),
TO_SIGNED(647,11),
TO_SIGNED(669,11),
TO_SIGNED(689,11),
TO_SIGNED(706,11),
TO_SIGNED(721,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(720,11),
TO_SIGNED(705,11),
TO_SIGNED(688,11),
TO_SIGNED(668,11),
TO_SIGNED(645,11),
TO_SIGNED(620,11),
TO_SIGNED(592,11),
TO_SIGNED(562,11),
TO_SIGNED(530,11),
TO_SIGNED(496,11),
TO_SIGNED(460,11),
TO_SIGNED(422,11),
TO_SIGNED(382,11),
TO_SIGNED(341,11),
TO_SIGNED(298,11),
TO_SIGNED(255,11),
TO_SIGNED(210,11),
TO_SIGNED(164,11),
TO_SIGNED(118,11),
TO_SIGNED(71,11),
TO_SIGNED(25,11),
TO_SIGNED(-22,11),
TO_SIGNED(-69,11),
TO_SIGNED(-116,11),
TO_SIGNED(-162,11),
TO_SIGNED(-208,11),
TO_SIGNED(-252,11),
TO_SIGNED(-296,11),
TO_SIGNED(-339,11),
TO_SIGNED(-380,11),
TO_SIGNED(-420,11),
TO_SIGNED(-458,11),
TO_SIGNED(-494,11),
TO_SIGNED(-529,11),
TO_SIGNED(-561,11),
TO_SIGNED(-591,11),
TO_SIGNED(-619,11),
TO_SIGNED(-644,11),
TO_SIGNED(-667,11),
TO_SIGNED(-687,11),
TO_SIGNED(-705,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-733,11),
TO_SIGNED(-721,11),
TO_SIGNED(-707,11),
TO_SIGNED(-690,11),
TO_SIGNED(-670,11),
TO_SIGNED(-648,11),
TO_SIGNED(-623,11),
TO_SIGNED(-596,11),
TO_SIGNED(-566,11),
TO_SIGNED(-534,11),
TO_SIGNED(-500,11),
TO_SIGNED(-464,11),
TO_SIGNED(-426,11),
TO_SIGNED(-387,11),
TO_SIGNED(-345,11),
TO_SIGNED(-303,11),
TO_SIGNED(-260,11),
TO_SIGNED(-215,11),
TO_SIGNED(-169,11),
TO_SIGNED(-123,11),
TO_SIGNED(-77,11),
TO_SIGNED(-30,11),
TO_SIGNED(17,11),
TO_SIGNED(64,11),
TO_SIGNED(111,11),
TO_SIGNED(157,11),
TO_SIGNED(203,11),
TO_SIGNED(247,11),
TO_SIGNED(291,11),
TO_SIGNED(334,11),
TO_SIGNED(375,11),
TO_SIGNED(415,11),
TO_SIGNED(454,11),
TO_SIGNED(490,11),
TO_SIGNED(525,11),
TO_SIGNED(557,11),
TO_SIGNED(588,11),
TO_SIGNED(616,11),
TO_SIGNED(641,11),
TO_SIGNED(664,11),
TO_SIGNED(685,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(709,11),
TO_SIGNED(692,11),
TO_SIGNED(673,11),
TO_SIGNED(651,11),
TO_SIGNED(626,11),
TO_SIGNED(599,11),
TO_SIGNED(569,11),
TO_SIGNED(538,11),
TO_SIGNED(504,11),
TO_SIGNED(468,11),
TO_SIGNED(430,11),
TO_SIGNED(391,11),
TO_SIGNED(350,11),
TO_SIGNED(308,11),
TO_SIGNED(265,11),
TO_SIGNED(220,11),
TO_SIGNED(175,11),
TO_SIGNED(129,11),
TO_SIGNED(82,11),
TO_SIGNED(35,11),
TO_SIGNED(-12,11),
TO_SIGNED(-59,11),
TO_SIGNED(-105,11),
TO_SIGNED(-152,11),
TO_SIGNED(-197,11),
TO_SIGNED(-242,11),
TO_SIGNED(-286,11),
TO_SIGNED(-329,11),
TO_SIGNED(-371,11),
TO_SIGNED(-411,11),
TO_SIGNED(-449,11),
TO_SIGNED(-486,11),
TO_SIGNED(-521,11),
TO_SIGNED(-554,11),
TO_SIGNED(-584,11),
TO_SIGNED(-613,11),
TO_SIGNED(-639,11),
TO_SIGNED(-662,11),
TO_SIGNED(-683,11),
TO_SIGNED(-701,11),
TO_SIGNED(-716,11),
TO_SIGNED(-729,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-711,11),
TO_SIGNED(-694,11),
TO_SIGNED(-675,11),
TO_SIGNED(-653,11),
TO_SIGNED(-629,11),
TO_SIGNED(-602,11),
TO_SIGNED(-573,11),
TO_SIGNED(-541,11),
TO_SIGNED(-508,11),
TO_SIGNED(-472,11),
TO_SIGNED(-435,11),
TO_SIGNED(-396,11),
TO_SIGNED(-355,11),
TO_SIGNED(-313,11),
TO_SIGNED(-270,11),
TO_SIGNED(-225,11),
TO_SIGNED(-180,11),
TO_SIGNED(-134,11),
TO_SIGNED(-87,11),
TO_SIGNED(-41,11),
TO_SIGNED(6,11),
TO_SIGNED(53,11),
TO_SIGNED(100,11),
TO_SIGNED(147,11),
TO_SIGNED(192,11),
TO_SIGNED(237,11),
TO_SIGNED(281,11),
TO_SIGNED(324,11),
TO_SIGNED(366,11),
TO_SIGNED(406,11),
TO_SIGNED(445,11),
TO_SIGNED(482,11),
TO_SIGNED(517,11),
TO_SIGNED(550,11),
TO_SIGNED(581,11),
TO_SIGNED(610,11),
TO_SIGNED(636,11),
TO_SIGNED(659,11),
TO_SIGNED(681,11),
TO_SIGNED(699,11),
TO_SIGNED(715,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(712,11),
TO_SIGNED(696,11),
TO_SIGNED(677,11),
TO_SIGNED(656,11),
TO_SIGNED(632,11),
TO_SIGNED(605,11),
TO_SIGNED(576,11),
TO_SIGNED(545,11),
TO_SIGNED(512,11),
TO_SIGNED(476,11),
TO_SIGNED(439,11),
TO_SIGNED(400,11),
TO_SIGNED(360,11),
TO_SIGNED(318,11),
TO_SIGNED(275,11),
TO_SIGNED(230,11),
TO_SIGNED(185,11),
TO_SIGNED(139,11),
TO_SIGNED(93,11),
TO_SIGNED(46,11),
TO_SIGNED(-1,11),
TO_SIGNED(-48,11),
TO_SIGNED(-95,11),
TO_SIGNED(-141,11),
TO_SIGNED(-187,11),
TO_SIGNED(-232,11),
TO_SIGNED(-276,11),
TO_SIGNED(-320,11),
TO_SIGNED(-362,11),
TO_SIGNED(-402,11),
TO_SIGNED(-441,11),
TO_SIGNED(-478,11),
TO_SIGNED(-513,11),
TO_SIGNED(-547,11),
TO_SIGNED(-578,11),
TO_SIGNED(-606,11),
TO_SIGNED(-633,11),
TO_SIGNED(-657,11),
TO_SIGNED(-678,11),
TO_SIGNED(-697,11),
TO_SIGNED(-713,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-714,11),
TO_SIGNED(-698,11),
TO_SIGNED(-680,11),
TO_SIGNED(-658,11),
TO_SIGNED(-635,11),
TO_SIGNED(-608,11),
TO_SIGNED(-580,11),
TO_SIGNED(-549,11),
TO_SIGNED(-516,11),
TO_SIGNED(-480,11),
TO_SIGNED(-443,11),
TO_SIGNED(-405,11),
TO_SIGNED(-364,11),
TO_SIGNED(-323,11),
TO_SIGNED(-279,11),
TO_SIGNED(-235,11),
TO_SIGNED(-190,11),
TO_SIGNED(-144,11),
TO_SIGNED(-98,11),
TO_SIGNED(-51,11),
TO_SIGNED(-4,11),
TO_SIGNED(43,11),
TO_SIGNED(90,11),
TO_SIGNED(136,11),
TO_SIGNED(182,11),
TO_SIGNED(227,11),
TO_SIGNED(272,11),
TO_SIGNED(315,11),
TO_SIGNED(357,11),
TO_SIGNED(397,11),
TO_SIGNED(437,11),
TO_SIGNED(474,11),
TO_SIGNED(509,11),
TO_SIGNED(543,11),
TO_SIGNED(574,11),
TO_SIGNED(603,11),
TO_SIGNED(630,11),
TO_SIGNED(654,11),
TO_SIGNED(676,11),
TO_SIGNED(695,11),
TO_SIGNED(711,11),
TO_SIGNED(725,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(716,11),
TO_SIGNED(700,11),
TO_SIGNED(682,11),
TO_SIGNED(661,11),
TO_SIGNED(637,11),
TO_SIGNED(611,11),
TO_SIGNED(583,11),
TO_SIGNED(552,11),
TO_SIGNED(519,11),
TO_SIGNED(485,11),
TO_SIGNED(448,11),
TO_SIGNED(409,11),
TO_SIGNED(369,11),
TO_SIGNED(327,11),
TO_SIGNED(284,11),
TO_SIGNED(240,11),
TO_SIGNED(195,11),
TO_SIGNED(150,11),
TO_SIGNED(103,11),
TO_SIGNED(57,11),
TO_SIGNED(10,11),
TO_SIGNED(-37,11),
TO_SIGNED(-84,11),
TO_SIGNED(-131,11),
TO_SIGNED(-177,11),
TO_SIGNED(-222,11),
TO_SIGNED(-267,11),
TO_SIGNED(-310,11),
TO_SIGNED(-352,11),
TO_SIGNED(-393,11),
TO_SIGNED(-432,11),
TO_SIGNED(-470,11),
TO_SIGNED(-505,11),
TO_SIGNED(-539,11),
TO_SIGNED(-571,11),
TO_SIGNED(-600,11),
TO_SIGNED(-627,11),
TO_SIGNED(-652,11),
TO_SIGNED(-674,11),
TO_SIGNED(-693,11),
TO_SIGNED(-710,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-702,11),
TO_SIGNED(-684,11),
TO_SIGNED(-663,11),
TO_SIGNED(-640,11),
TO_SIGNED(-615,11),
TO_SIGNED(-586,11),
TO_SIGNED(-556,11),
TO_SIGNED(-523,11),
TO_SIGNED(-489,11),
TO_SIGNED(-452,11),
TO_SIGNED(-414,11),
TO_SIGNED(-374,11),
TO_SIGNED(-332,11),
TO_SIGNED(-289,11),
TO_SIGNED(-245,11),
TO_SIGNED(-201,11),
TO_SIGNED(-155,11),
TO_SIGNED(-109,11),
TO_SIGNED(-62,11),
TO_SIGNED(-15,11),
TO_SIGNED(32,11),
TO_SIGNED(79,11),
TO_SIGNED(125,11),
TO_SIGNED(172,11),
TO_SIGNED(217,11),
TO_SIGNED(262,11),
TO_SIGNED(305,11),
TO_SIGNED(347,11),
TO_SIGNED(388,11),
TO_SIGNED(428,11),
TO_SIGNED(466,11),
TO_SIGNED(501,11),
TO_SIGNED(535,11),
TO_SIGNED(567,11),
TO_SIGNED(597,11),
TO_SIGNED(624,11),
TO_SIGNED(649,11),
TO_SIGNED(671,11),
TO_SIGNED(691,11),
TO_SIGNED(708,11),
TO_SIGNED(722,11),
TO_SIGNED(733,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(704,11),
TO_SIGNED(686,11),
TO_SIGNED(666,11),
TO_SIGNED(643,11),
TO_SIGNED(618,11),
TO_SIGNED(590,11),
TO_SIGNED(559,11),
TO_SIGNED(527,11),
TO_SIGNED(493,11),
TO_SIGNED(456,11),
TO_SIGNED(418,11),
TO_SIGNED(378,11),
TO_SIGNED(337,11),
TO_SIGNED(294,11),
TO_SIGNED(250,11),
TO_SIGNED(206,11),
TO_SIGNED(160,11),
TO_SIGNED(114,11),
TO_SIGNED(67,11),
TO_SIGNED(20,11),
TO_SIGNED(-27,11),
TO_SIGNED(-74,11),
TO_SIGNED(-120,11),
TO_SIGNED(-166,11),
TO_SIGNED(-212,11),
TO_SIGNED(-257,11),
TO_SIGNED(-300,11),
TO_SIGNED(-343,11),
TO_SIGNED(-384,11),
TO_SIGNED(-423,11),
TO_SIGNED(-461,11),
TO_SIGNED(-497,11),
TO_SIGNED(-532,11),
TO_SIGNED(-564,11),
TO_SIGNED(-594,11),
TO_SIGNED(-621,11),
TO_SIGNED(-646,11),
TO_SIGNED(-669,11),
TO_SIGNED(-689,11),
TO_SIGNED(-706,11),
TO_SIGNED(-721,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-720,11),
TO_SIGNED(-706,11),
TO_SIGNED(-688,11),
TO_SIGNED(-668,11),
TO_SIGNED(-646,11),
TO_SIGNED(-621,11),
TO_SIGNED(-593,11),
TO_SIGNED(-563,11),
TO_SIGNED(-531,11),
TO_SIGNED(-497,11),
TO_SIGNED(-460,11),
TO_SIGNED(-422,11),
TO_SIGNED(-383,11),
TO_SIGNED(-342,11),
TO_SIGNED(-299,11),
TO_SIGNED(-256,11),
TO_SIGNED(-211,11),
TO_SIGNED(-165,11),
TO_SIGNED(-119,11),
TO_SIGNED(-73,11),
TO_SIGNED(-26,11),
TO_SIGNED(21,11),
TO_SIGNED(68,11),
TO_SIGNED(115,11),
TO_SIGNED(161,11),
TO_SIGNED(207,11),
TO_SIGNED(251,11),
TO_SIGNED(295,11),
TO_SIGNED(338,11),
TO_SIGNED(379,11),
TO_SIGNED(419,11),
TO_SIGNED(457,11),
TO_SIGNED(493,11),
TO_SIGNED(528,11),
TO_SIGNED(560,11),
TO_SIGNED(590,11),
TO_SIGNED(618,11),
TO_SIGNED(644,11),
TO_SIGNED(666,11),
TO_SIGNED(687,11),
TO_SIGNED(704,11),
TO_SIGNED(719,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(671,11),
TO_SIGNED(648,11),
TO_SIGNED(624,11),
TO_SIGNED(596,11),
TO_SIGNED(567,11),
TO_SIGNED(535,11),
TO_SIGNED(501,11),
TO_SIGNED(465,11),
TO_SIGNED(427,11),
TO_SIGNED(387,11),
TO_SIGNED(346,11),
TO_SIGNED(304,11),
TO_SIGNED(261,11),
TO_SIGNED(216,11),
TO_SIGNED(171,11),
TO_SIGNED(124,11),
TO_SIGNED(78,11),
TO_SIGNED(31,11),
TO_SIGNED(-16,11),
TO_SIGNED(-63,11),
TO_SIGNED(-110,11),
TO_SIGNED(-156,11),
TO_SIGNED(-202,11),
TO_SIGNED(-246,11),
TO_SIGNED(-290,11),
TO_SIGNED(-333,11),
TO_SIGNED(-375,11),
TO_SIGNED(-415,11),
TO_SIGNED(-453,11),
TO_SIGNED(-489,11),
TO_SIGNED(-524,11),
TO_SIGNED(-557,11),
TO_SIGNED(-587,11),
TO_SIGNED(-615,11),
TO_SIGNED(-641,11),
TO_SIGNED(-664,11),
TO_SIGNED(-685,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-730,11),
TO_SIGNED(-739,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-693,11),
TO_SIGNED(-673,11),
TO_SIGNED(-651,11),
TO_SIGNED(-627,11),
TO_SIGNED(-599,11),
TO_SIGNED(-570,11),
TO_SIGNED(-538,11),
TO_SIGNED(-505,11),
TO_SIGNED(-469,11),
TO_SIGNED(-431,11),
TO_SIGNED(-392,11),
TO_SIGNED(-351,11),
TO_SIGNED(-309,11),
TO_SIGNED(-266,11),
TO_SIGNED(-221,11),
TO_SIGNED(-176,11),
TO_SIGNED(-130,11),
TO_SIGNED(-83,11),
TO_SIGNED(-36,11),
TO_SIGNED(11,11),
TO_SIGNED(58,11),
TO_SIGNED(104,11),
TO_SIGNED(151,11),
TO_SIGNED(196,11),
TO_SIGNED(241,11),
TO_SIGNED(285,11),
TO_SIGNED(328,11),
TO_SIGNED(370,11),
TO_SIGNED(410,11),
TO_SIGNED(449,11),
TO_SIGNED(485,11),
TO_SIGNED(520,11),
TO_SIGNED(553,11),
TO_SIGNED(584,11),
TO_SIGNED(612,11),
TO_SIGNED(638,11),
TO_SIGNED(661,11),
TO_SIGNED(682,11),
TO_SIGNED(700,11),
TO_SIGNED(716,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(725,11),
TO_SIGNED(711,11),
TO_SIGNED(695,11),
TO_SIGNED(675,11),
TO_SIGNED(654,11),
TO_SIGNED(629,11),
TO_SIGNED(603,11),
TO_SIGNED(574,11),
TO_SIGNED(542,11),
TO_SIGNED(509,11),
TO_SIGNED(473,11),
TO_SIGNED(436,11),
TO_SIGNED(397,11),
TO_SIGNED(356,11),
TO_SIGNED(314,11),
TO_SIGNED(271,11),
TO_SIGNED(226,11),
TO_SIGNED(181,11),
TO_SIGNED(135,11),
TO_SIGNED(88,11),
TO_SIGNED(42,11),
TO_SIGNED(-5,11),
TO_SIGNED(-52,11),
TO_SIGNED(-99,11),
TO_SIGNED(-145,11),
TO_SIGNED(-191,11),
TO_SIGNED(-236,11),
TO_SIGNED(-280,11),
TO_SIGNED(-323,11),
TO_SIGNED(-365,11),
TO_SIGNED(-406,11),
TO_SIGNED(-444,11),
TO_SIGNED(-481,11),
TO_SIGNED(-516,11),
TO_SIGNED(-549,11),
TO_SIGNED(-580,11),
TO_SIGNED(-609,11),
TO_SIGNED(-635,11),
TO_SIGNED(-659,11),
TO_SIGNED(-680,11),
TO_SIGNED(-699,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-736,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-678,11),
TO_SIGNED(-656,11),
TO_SIGNED(-632,11),
TO_SIGNED(-606,11),
TO_SIGNED(-577,11),
TO_SIGNED(-546,11),
TO_SIGNED(-512,11),
TO_SIGNED(-477,11),
TO_SIGNED(-440,11),
TO_SIGNED(-401,11),
TO_SIGNED(-361,11),
TO_SIGNED(-319,11),
TO_SIGNED(-275,11),
TO_SIGNED(-231,11),
TO_SIGNED(-186,11),
TO_SIGNED(-140,11),
TO_SIGNED(-94,11),
TO_SIGNED(-47,11),
TO_SIGNED(0,11),
TO_SIGNED(47,11),
TO_SIGNED(94,11),
TO_SIGNED(140,11),
TO_SIGNED(186,11),
TO_SIGNED(231,11),
TO_SIGNED(275,11),
TO_SIGNED(319,11),
TO_SIGNED(361,11),
TO_SIGNED(401,11),
TO_SIGNED(440,11),
TO_SIGNED(477,11),
TO_SIGNED(512,11),
TO_SIGNED(546,11),
TO_SIGNED(577,11),
TO_SIGNED(606,11),
TO_SIGNED(632,11),
TO_SIGNED(656,11),
TO_SIGNED(678,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(736,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(699,11),
TO_SIGNED(680,11),
TO_SIGNED(659,11),
TO_SIGNED(635,11),
TO_SIGNED(609,11),
TO_SIGNED(580,11),
TO_SIGNED(549,11),
TO_SIGNED(516,11),
TO_SIGNED(481,11),
TO_SIGNED(444,11),
TO_SIGNED(406,11),
TO_SIGNED(365,11),
TO_SIGNED(323,11),
TO_SIGNED(280,11),
TO_SIGNED(236,11),
TO_SIGNED(191,11),
TO_SIGNED(145,11),
TO_SIGNED(99,11),
TO_SIGNED(52,11),
TO_SIGNED(5,11),
TO_SIGNED(-42,11),
TO_SIGNED(-88,11),
TO_SIGNED(-135,11),
TO_SIGNED(-181,11),
TO_SIGNED(-226,11),
TO_SIGNED(-271,11),
TO_SIGNED(-314,11),
TO_SIGNED(-356,11),
TO_SIGNED(-397,11),
TO_SIGNED(-436,11),
TO_SIGNED(-473,11),
TO_SIGNED(-509,11),
TO_SIGNED(-542,11),
TO_SIGNED(-574,11),
TO_SIGNED(-603,11),
TO_SIGNED(-629,11),
TO_SIGNED(-654,11),
TO_SIGNED(-675,11),
TO_SIGNED(-695,11),
TO_SIGNED(-711,11),
TO_SIGNED(-725,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-716,11),
TO_SIGNED(-700,11),
TO_SIGNED(-682,11),
TO_SIGNED(-661,11),
TO_SIGNED(-638,11),
TO_SIGNED(-612,11),
TO_SIGNED(-584,11),
TO_SIGNED(-553,11),
TO_SIGNED(-520,11),
TO_SIGNED(-485,11),
TO_SIGNED(-449,11),
TO_SIGNED(-410,11),
TO_SIGNED(-370,11),
TO_SIGNED(-328,11),
TO_SIGNED(-285,11),
TO_SIGNED(-241,11),
TO_SIGNED(-196,11),
TO_SIGNED(-151,11),
TO_SIGNED(-104,11),
TO_SIGNED(-58,11),
TO_SIGNED(-11,11),
TO_SIGNED(36,11),
TO_SIGNED(83,11),
TO_SIGNED(130,11),
TO_SIGNED(176,11),
TO_SIGNED(221,11),
TO_SIGNED(266,11),
TO_SIGNED(309,11),
TO_SIGNED(351,11),
TO_SIGNED(392,11),
TO_SIGNED(431,11),
TO_SIGNED(469,11),
TO_SIGNED(505,11),
TO_SIGNED(538,11),
TO_SIGNED(570,11),
TO_SIGNED(599,11),
TO_SIGNED(627,11),
TO_SIGNED(651,11),
TO_SIGNED(673,11),
TO_SIGNED(693,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(739,11),
TO_SIGNED(730,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(685,11),
TO_SIGNED(664,11),
TO_SIGNED(641,11),
TO_SIGNED(615,11),
TO_SIGNED(587,11),
TO_SIGNED(557,11),
TO_SIGNED(524,11),
TO_SIGNED(489,11),
TO_SIGNED(453,11),
TO_SIGNED(415,11),
TO_SIGNED(375,11),
TO_SIGNED(333,11),
TO_SIGNED(290,11),
TO_SIGNED(246,11),
TO_SIGNED(202,11),
TO_SIGNED(156,11),
TO_SIGNED(110,11),
TO_SIGNED(63,11),
TO_SIGNED(16,11),
TO_SIGNED(-31,11),
TO_SIGNED(-78,11),
TO_SIGNED(-124,11),
TO_SIGNED(-171,11),
TO_SIGNED(-216,11),
TO_SIGNED(-261,11),
TO_SIGNED(-304,11),
TO_SIGNED(-346,11),
TO_SIGNED(-387,11),
TO_SIGNED(-427,11),
TO_SIGNED(-465,11),
TO_SIGNED(-501,11),
TO_SIGNED(-535,11),
TO_SIGNED(-567,11),
TO_SIGNED(-596,11),
TO_SIGNED(-624,11),
TO_SIGNED(-648,11),
TO_SIGNED(-671,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-719,11),
TO_SIGNED(-704,11),
TO_SIGNED(-687,11),
TO_SIGNED(-666,11),
TO_SIGNED(-644,11),
TO_SIGNED(-618,11),
TO_SIGNED(-590,11),
TO_SIGNED(-560,11),
TO_SIGNED(-528,11),
TO_SIGNED(-493,11),
TO_SIGNED(-457,11),
TO_SIGNED(-419,11),
TO_SIGNED(-379,11),
TO_SIGNED(-338,11),
TO_SIGNED(-295,11),
TO_SIGNED(-251,11),
TO_SIGNED(-207,11),
TO_SIGNED(-161,11),
TO_SIGNED(-115,11),
TO_SIGNED(-68,11),
TO_SIGNED(-21,11),
TO_SIGNED(26,11),
TO_SIGNED(73,11),
TO_SIGNED(119,11),
TO_SIGNED(165,11),
TO_SIGNED(211,11),
TO_SIGNED(256,11),
TO_SIGNED(299,11),
TO_SIGNED(342,11),
TO_SIGNED(383,11),
TO_SIGNED(422,11),
TO_SIGNED(460,11),
TO_SIGNED(497,11),
TO_SIGNED(531,11),
TO_SIGNED(563,11),
TO_SIGNED(593,11),
TO_SIGNED(621,11),
TO_SIGNED(646,11),
TO_SIGNED(668,11),
TO_SIGNED(688,11),
TO_SIGNED(706,11),
TO_SIGNED(720,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(721,11),
TO_SIGNED(706,11),
TO_SIGNED(689,11),
TO_SIGNED(669,11),
TO_SIGNED(646,11),
TO_SIGNED(621,11),
TO_SIGNED(594,11),
TO_SIGNED(564,11),
TO_SIGNED(532,11),
TO_SIGNED(497,11),
TO_SIGNED(461,11),
TO_SIGNED(423,11),
TO_SIGNED(384,11),
TO_SIGNED(343,11),
TO_SIGNED(300,11),
TO_SIGNED(257,11),
TO_SIGNED(212,11),
TO_SIGNED(166,11),
TO_SIGNED(120,11),
TO_SIGNED(74,11),
TO_SIGNED(27,11),
TO_SIGNED(-20,11),
TO_SIGNED(-67,11),
TO_SIGNED(-114,11),
TO_SIGNED(-160,11),
TO_SIGNED(-206,11),
TO_SIGNED(-250,11),
TO_SIGNED(-294,11),
TO_SIGNED(-337,11),
TO_SIGNED(-378,11),
TO_SIGNED(-418,11),
TO_SIGNED(-456,11),
TO_SIGNED(-493,11),
TO_SIGNED(-527,11),
TO_SIGNED(-559,11),
TO_SIGNED(-590,11),
TO_SIGNED(-618,11),
TO_SIGNED(-643,11),
TO_SIGNED(-666,11),
TO_SIGNED(-686,11),
TO_SIGNED(-704,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-733,11),
TO_SIGNED(-722,11),
TO_SIGNED(-708,11),
TO_SIGNED(-691,11),
TO_SIGNED(-671,11),
TO_SIGNED(-649,11),
TO_SIGNED(-624,11),
TO_SIGNED(-597,11),
TO_SIGNED(-567,11),
TO_SIGNED(-535,11),
TO_SIGNED(-501,11),
TO_SIGNED(-466,11),
TO_SIGNED(-428,11),
TO_SIGNED(-388,11),
TO_SIGNED(-347,11),
TO_SIGNED(-305,11),
TO_SIGNED(-262,11),
TO_SIGNED(-217,11),
TO_SIGNED(-172,11),
TO_SIGNED(-125,11),
TO_SIGNED(-79,11),
TO_SIGNED(-32,11),
TO_SIGNED(15,11),
TO_SIGNED(62,11),
TO_SIGNED(109,11),
TO_SIGNED(155,11),
TO_SIGNED(201,11),
TO_SIGNED(245,11),
TO_SIGNED(289,11),
TO_SIGNED(332,11),
TO_SIGNED(374,11),
TO_SIGNED(414,11),
TO_SIGNED(452,11),
TO_SIGNED(489,11),
TO_SIGNED(523,11),
TO_SIGNED(556,11),
TO_SIGNED(586,11),
TO_SIGNED(615,11),
TO_SIGNED(640,11),
TO_SIGNED(663,11),
TO_SIGNED(684,11),
TO_SIGNED(702,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(710,11),
TO_SIGNED(693,11),
TO_SIGNED(674,11),
TO_SIGNED(652,11),
TO_SIGNED(627,11),
TO_SIGNED(600,11),
TO_SIGNED(571,11),
TO_SIGNED(539,11),
TO_SIGNED(505,11),
TO_SIGNED(470,11),
TO_SIGNED(432,11),
TO_SIGNED(393,11),
TO_SIGNED(352,11),
TO_SIGNED(310,11),
TO_SIGNED(267,11),
TO_SIGNED(222,11),
TO_SIGNED(177,11),
TO_SIGNED(131,11),
TO_SIGNED(84,11),
TO_SIGNED(37,11),
TO_SIGNED(-10,11),
TO_SIGNED(-57,11),
TO_SIGNED(-103,11),
TO_SIGNED(-150,11),
TO_SIGNED(-195,11),
TO_SIGNED(-240,11),
TO_SIGNED(-284,11),
TO_SIGNED(-327,11),
TO_SIGNED(-369,11),
TO_SIGNED(-409,11),
TO_SIGNED(-448,11),
TO_SIGNED(-485,11),
TO_SIGNED(-519,11),
TO_SIGNED(-552,11),
TO_SIGNED(-583,11),
TO_SIGNED(-611,11),
TO_SIGNED(-637,11),
TO_SIGNED(-661,11),
TO_SIGNED(-682,11),
TO_SIGNED(-700,11),
TO_SIGNED(-716,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-725,11),
TO_SIGNED(-711,11),
TO_SIGNED(-695,11),
TO_SIGNED(-676,11),
TO_SIGNED(-654,11),
TO_SIGNED(-630,11),
TO_SIGNED(-603,11),
TO_SIGNED(-574,11),
TO_SIGNED(-543,11),
TO_SIGNED(-509,11),
TO_SIGNED(-474,11),
TO_SIGNED(-437,11),
TO_SIGNED(-397,11),
TO_SIGNED(-357,11),
TO_SIGNED(-315,11),
TO_SIGNED(-272,11),
TO_SIGNED(-227,11),
TO_SIGNED(-182,11),
TO_SIGNED(-136,11),
TO_SIGNED(-90,11),
TO_SIGNED(-43,11),
TO_SIGNED(4,11),
TO_SIGNED(51,11),
TO_SIGNED(98,11),
TO_SIGNED(144,11),
TO_SIGNED(190,11),
TO_SIGNED(235,11),
TO_SIGNED(279,11),
TO_SIGNED(323,11),
TO_SIGNED(364,11),
TO_SIGNED(405,11),
TO_SIGNED(443,11),
TO_SIGNED(480,11),
TO_SIGNED(516,11),
TO_SIGNED(549,11),
TO_SIGNED(580,11),
TO_SIGNED(608,11),
TO_SIGNED(635,11),
TO_SIGNED(658,11),
TO_SIGNED(680,11),
TO_SIGNED(698,11),
TO_SIGNED(714,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(713,11),
TO_SIGNED(697,11),
TO_SIGNED(678,11),
TO_SIGNED(657,11),
TO_SIGNED(633,11),
TO_SIGNED(606,11),
TO_SIGNED(578,11),
TO_SIGNED(547,11),
TO_SIGNED(513,11),
TO_SIGNED(478,11),
TO_SIGNED(441,11),
TO_SIGNED(402,11),
TO_SIGNED(362,11),
TO_SIGNED(320,11),
TO_SIGNED(276,11),
TO_SIGNED(232,11),
TO_SIGNED(187,11),
TO_SIGNED(141,11),
TO_SIGNED(95,11),
TO_SIGNED(48,11),
TO_SIGNED(1,11),
TO_SIGNED(-46,11),
TO_SIGNED(-93,11),
TO_SIGNED(-139,11),
TO_SIGNED(-185,11),
TO_SIGNED(-230,11),
TO_SIGNED(-275,11),
TO_SIGNED(-318,11),
TO_SIGNED(-360,11),
TO_SIGNED(-400,11),
TO_SIGNED(-439,11),
TO_SIGNED(-476,11),
TO_SIGNED(-512,11),
TO_SIGNED(-545,11),
TO_SIGNED(-576,11),
TO_SIGNED(-605,11),
TO_SIGNED(-632,11),
TO_SIGNED(-656,11),
TO_SIGNED(-677,11),
TO_SIGNED(-696,11),
TO_SIGNED(-712,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-715,11),
TO_SIGNED(-699,11),
TO_SIGNED(-681,11),
TO_SIGNED(-659,11),
TO_SIGNED(-636,11),
TO_SIGNED(-610,11),
TO_SIGNED(-581,11),
TO_SIGNED(-550,11),
TO_SIGNED(-517,11),
TO_SIGNED(-482,11),
TO_SIGNED(-445,11),
TO_SIGNED(-406,11),
TO_SIGNED(-366,11),
TO_SIGNED(-324,11),
TO_SIGNED(-281,11),
TO_SIGNED(-237,11),
TO_SIGNED(-192,11),
TO_SIGNED(-147,11),
TO_SIGNED(-100,11),
TO_SIGNED(-53,11),
TO_SIGNED(-6,11),
TO_SIGNED(41,11),
TO_SIGNED(87,11),
TO_SIGNED(134,11),
TO_SIGNED(180,11),
TO_SIGNED(225,11),
TO_SIGNED(270,11),
TO_SIGNED(313,11),
TO_SIGNED(355,11),
TO_SIGNED(396,11),
TO_SIGNED(435,11),
TO_SIGNED(472,11),
TO_SIGNED(508,11),
TO_SIGNED(541,11),
TO_SIGNED(573,11),
TO_SIGNED(602,11),
TO_SIGNED(629,11),
TO_SIGNED(653,11),
TO_SIGNED(675,11),
TO_SIGNED(694,11),
TO_SIGNED(711,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(729,11),
TO_SIGNED(716,11),
TO_SIGNED(701,11),
TO_SIGNED(683,11),
TO_SIGNED(662,11),
TO_SIGNED(639,11),
TO_SIGNED(613,11),
TO_SIGNED(584,11),
TO_SIGNED(554,11),
TO_SIGNED(521,11),
TO_SIGNED(486,11),
TO_SIGNED(449,11),
TO_SIGNED(411,11),
TO_SIGNED(371,11),
TO_SIGNED(329,11),
TO_SIGNED(286,11),
TO_SIGNED(242,11),
TO_SIGNED(197,11),
TO_SIGNED(152,11),
TO_SIGNED(105,11),
TO_SIGNED(59,11),
TO_SIGNED(12,11),
TO_SIGNED(-35,11),
TO_SIGNED(-82,11),
TO_SIGNED(-129,11),
TO_SIGNED(-175,11),
TO_SIGNED(-220,11),
TO_SIGNED(-265,11),
TO_SIGNED(-308,11),
TO_SIGNED(-350,11),
TO_SIGNED(-391,11),
TO_SIGNED(-430,11),
TO_SIGNED(-468,11),
TO_SIGNED(-504,11),
TO_SIGNED(-538,11),
TO_SIGNED(-569,11),
TO_SIGNED(-599,11),
TO_SIGNED(-626,11),
TO_SIGNED(-651,11),
TO_SIGNED(-673,11),
TO_SIGNED(-692,11),
TO_SIGNED(-709,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-685,11),
TO_SIGNED(-664,11),
TO_SIGNED(-641,11),
TO_SIGNED(-616,11),
TO_SIGNED(-588,11),
TO_SIGNED(-557,11),
TO_SIGNED(-525,11),
TO_SIGNED(-490,11),
TO_SIGNED(-454,11),
TO_SIGNED(-415,11),
TO_SIGNED(-375,11),
TO_SIGNED(-334,11),
TO_SIGNED(-291,11),
TO_SIGNED(-247,11),
TO_SIGNED(-203,11),
TO_SIGNED(-157,11),
TO_SIGNED(-111,11),
TO_SIGNED(-64,11),
TO_SIGNED(-17,11),
TO_SIGNED(30,11),
TO_SIGNED(77,11),
TO_SIGNED(123,11),
TO_SIGNED(169,11),
TO_SIGNED(215,11),
TO_SIGNED(260,11),
TO_SIGNED(303,11),
TO_SIGNED(345,11),
TO_SIGNED(387,11),
TO_SIGNED(426,11),
TO_SIGNED(464,11),
TO_SIGNED(500,11),
TO_SIGNED(534,11),
TO_SIGNED(566,11),
TO_SIGNED(596,11),
TO_SIGNED(623,11),
TO_SIGNED(648,11),
TO_SIGNED(670,11),
TO_SIGNED(690,11),
TO_SIGNED(707,11),
TO_SIGNED(721,11),
TO_SIGNED(733,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(705,11),
TO_SIGNED(687,11),
TO_SIGNED(667,11),
TO_SIGNED(644,11),
TO_SIGNED(619,11),
TO_SIGNED(591,11),
TO_SIGNED(561,11),
TO_SIGNED(529,11),
TO_SIGNED(494,11),
TO_SIGNED(458,11),
TO_SIGNED(420,11),
TO_SIGNED(380,11),
TO_SIGNED(339,11),
TO_SIGNED(296,11),
TO_SIGNED(252,11),
TO_SIGNED(208,11),
TO_SIGNED(162,11),
TO_SIGNED(116,11),
TO_SIGNED(69,11),
TO_SIGNED(22,11),
TO_SIGNED(-25,11),
TO_SIGNED(-71,11),
TO_SIGNED(-118,11),
TO_SIGNED(-164,11),
TO_SIGNED(-210,11),
TO_SIGNED(-255,11),
TO_SIGNED(-298,11),
TO_SIGNED(-341,11),
TO_SIGNED(-382,11),
TO_SIGNED(-422,11),
TO_SIGNED(-460,11),
TO_SIGNED(-496,11),
TO_SIGNED(-530,11),
TO_SIGNED(-562,11),
TO_SIGNED(-592,11),
TO_SIGNED(-620,11),
TO_SIGNED(-645,11),
TO_SIGNED(-668,11),
TO_SIGNED(-688,11),
TO_SIGNED(-705,11),
TO_SIGNED(-720,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-721,11),
TO_SIGNED(-706,11),
TO_SIGNED(-689,11),
TO_SIGNED(-669,11),
TO_SIGNED(-647,11),
TO_SIGNED(-622,11),
TO_SIGNED(-594,11),
TO_SIGNED(-564,11),
TO_SIGNED(-532,11),
TO_SIGNED(-498,11),
TO_SIGNED(-462,11),
TO_SIGNED(-424,11),
TO_SIGNED(-385,11),
TO_SIGNED(-344,11),
TO_SIGNED(-301,11),
TO_SIGNED(-258,11),
TO_SIGNED(-213,11),
TO_SIGNED(-167,11),
TO_SIGNED(-121,11),
TO_SIGNED(-75,11),
TO_SIGNED(-28,11),
TO_SIGNED(19,11),
TO_SIGNED(66,11),
TO_SIGNED(113,11),
TO_SIGNED(159,11),
TO_SIGNED(205,11),
TO_SIGNED(249,11),
TO_SIGNED(293,11),
TO_SIGNED(336,11),
TO_SIGNED(377,11),
TO_SIGNED(417,11),
TO_SIGNED(455,11),
TO_SIGNED(492,11),
TO_SIGNED(526,11),
TO_SIGNED(559,11),
TO_SIGNED(589,11),
TO_SIGNED(617,11),
TO_SIGNED(642,11),
TO_SIGNED(665,11),
TO_SIGNED(686,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(708,11),
TO_SIGNED(691,11),
TO_SIGNED(672,11),
TO_SIGNED(650,11),
TO_SIGNED(625,11),
TO_SIGNED(598,11),
TO_SIGNED(568,11),
TO_SIGNED(536,11),
TO_SIGNED(502,11),
TO_SIGNED(466,11),
TO_SIGNED(429,11),
TO_SIGNED(389,11),
TO_SIGNED(348,11),
TO_SIGNED(306,11),
TO_SIGNED(263,11),
TO_SIGNED(218,11),
TO_SIGNED(173,11),
TO_SIGNED(127,11),
TO_SIGNED(80,11),
TO_SIGNED(33,11),
TO_SIGNED(-14,11),
TO_SIGNED(-61,11),
TO_SIGNED(-108,11),
TO_SIGNED(-154,11),
TO_SIGNED(-200,11),
TO_SIGNED(-244,11),
TO_SIGNED(-288,11),
TO_SIGNED(-331,11),
TO_SIGNED(-373,11),
TO_SIGNED(-413,11),
TO_SIGNED(-451,11),
TO_SIGNED(-488,11),
TO_SIGNED(-523,11),
TO_SIGNED(-555,11),
TO_SIGNED(-586,11),
TO_SIGNED(-614,11),
TO_SIGNED(-640,11),
TO_SIGNED(-663,11),
TO_SIGNED(-684,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-729,11),
TO_SIGNED(-739,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-710,11),
TO_SIGNED(-693,11),
TO_SIGNED(-674,11),
TO_SIGNED(-652,11),
TO_SIGNED(-628,11),
TO_SIGNED(-601,11),
TO_SIGNED(-571,11),
TO_SIGNED(-540,11),
TO_SIGNED(-506,11),
TO_SIGNED(-471,11),
TO_SIGNED(-433,11),
TO_SIGNED(-394,11),
TO_SIGNED(-353,11),
TO_SIGNED(-311,11),
TO_SIGNED(-268,11),
TO_SIGNED(-223,11),
TO_SIGNED(-178,11),
TO_SIGNED(-132,11),
TO_SIGNED(-85,11),
TO_SIGNED(-38,11),
TO_SIGNED(9,11),
TO_SIGNED(56,11),
TO_SIGNED(102,11),
TO_SIGNED(149,11),
TO_SIGNED(194,11),
TO_SIGNED(239,11),
TO_SIGNED(283,11),
TO_SIGNED(326,11),
TO_SIGNED(368,11),
TO_SIGNED(408,11),
TO_SIGNED(447,11),
TO_SIGNED(484,11),
TO_SIGNED(519,11),
TO_SIGNED(552,11),
TO_SIGNED(582,11),
TO_SIGNED(611,11),
TO_SIGNED(637,11),
TO_SIGNED(660,11),
TO_SIGNED(681,11),
TO_SIGNED(700,11),
TO_SIGNED(715,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(736,11),
TO_SIGNED(725,11),
TO_SIGNED(712,11),
TO_SIGNED(695,11),
TO_SIGNED(676,11),
TO_SIGNED(655,11),
TO_SIGNED(631,11),
TO_SIGNED(604,11),
TO_SIGNED(575,11),
TO_SIGNED(544,11),
TO_SIGNED(510,11),
TO_SIGNED(475,11),
TO_SIGNED(437,11),
TO_SIGNED(398,11),
TO_SIGNED(358,11),
TO_SIGNED(316,11),
TO_SIGNED(273,11),
TO_SIGNED(228,11),
TO_SIGNED(183,11),
TO_SIGNED(137,11),
TO_SIGNED(91,11),
TO_SIGNED(44,11),
TO_SIGNED(-3,11),
TO_SIGNED(-50,11),
TO_SIGNED(-97,11),
TO_SIGNED(-143,11),
TO_SIGNED(-189,11),
TO_SIGNED(-234,11),
TO_SIGNED(-278,11),
TO_SIGNED(-322,11),
TO_SIGNED(-363,11),
TO_SIGNED(-404,11),
TO_SIGNED(-443,11),
TO_SIGNED(-480,11),
TO_SIGNED(-515,11),
TO_SIGNED(-548,11),
TO_SIGNED(-579,11),
TO_SIGNED(-608,11),
TO_SIGNED(-634,11),
TO_SIGNED(-658,11),
TO_SIGNED(-679,11),
TO_SIGNED(-698,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-679,11),
TO_SIGNED(-657,11),
TO_SIGNED(-633,11),
TO_SIGNED(-607,11),
TO_SIGNED(-578,11),
TO_SIGNED(-547,11),
TO_SIGNED(-514,11),
TO_SIGNED(-479,11),
TO_SIGNED(-442,11),
TO_SIGNED(-403,11),
TO_SIGNED(-362,11),
TO_SIGNED(-321,11),
TO_SIGNED(-277,11),
TO_SIGNED(-233,11),
TO_SIGNED(-188,11),
TO_SIGNED(-142,11),
TO_SIGNED(-96,11),
TO_SIGNED(-49,11),
TO_SIGNED(-2,11),
TO_SIGNED(45,11),
TO_SIGNED(92,11),
TO_SIGNED(138,11),
TO_SIGNED(184,11),
TO_SIGNED(229,11),
TO_SIGNED(274,11),
TO_SIGNED(317,11),
TO_SIGNED(359,11),
TO_SIGNED(399,11),
TO_SIGNED(438,11),
TO_SIGNED(476,11),
TO_SIGNED(511,11),
TO_SIGNED(544,11),
TO_SIGNED(576,11),
TO_SIGNED(605,11),
TO_SIGNED(631,11),
TO_SIGNED(655,11),
TO_SIGNED(677,11),
TO_SIGNED(696,11),
TO_SIGNED(712,11),
TO_SIGNED(725,11),
TO_SIGNED(736,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(715,11),
TO_SIGNED(699,11),
TO_SIGNED(681,11),
TO_SIGNED(660,11),
TO_SIGNED(636,11),
TO_SIGNED(610,11),
TO_SIGNED(582,11),
TO_SIGNED(551,11),
TO_SIGNED(518,11),
TO_SIGNED(483,11),
TO_SIGNED(446,11),
TO_SIGNED(407,11),
TO_SIGNED(367,11),
TO_SIGNED(325,11),
TO_SIGNED(282,11),
TO_SIGNED(238,11),
TO_SIGNED(193,11),
TO_SIGNED(148,11),
TO_SIGNED(101,11),
TO_SIGNED(54,11),
TO_SIGNED(7,11),
TO_SIGNED(-40,11),
TO_SIGNED(-86,11),
TO_SIGNED(-133,11),
TO_SIGNED(-179,11),
TO_SIGNED(-224,11),
TO_SIGNED(-269,11),
TO_SIGNED(-312,11),
TO_SIGNED(-354,11),
TO_SIGNED(-395,11),
TO_SIGNED(-434,11),
TO_SIGNED(-471,11),
TO_SIGNED(-507,11),
TO_SIGNED(-541,11),
TO_SIGNED(-572,11),
TO_SIGNED(-601,11),
TO_SIGNED(-628,11),
TO_SIGNED(-653,11),
TO_SIGNED(-675,11),
TO_SIGNED(-694,11),
TO_SIGNED(-710,11),
TO_SIGNED(-724,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-701,11),
TO_SIGNED(-683,11),
TO_SIGNED(-662,11),
TO_SIGNED(-639,11),
TO_SIGNED(-613,11),
TO_SIGNED(-585,11),
TO_SIGNED(-554,11),
TO_SIGNED(-522,11),
TO_SIGNED(-487,11),
TO_SIGNED(-450,11),
TO_SIGNED(-412,11),
TO_SIGNED(-372,11),
TO_SIGNED(-330,11),
TO_SIGNED(-287,11),
TO_SIGNED(-243,11),
TO_SIGNED(-198,11),
TO_SIGNED(-153,11),
TO_SIGNED(-106,11),
TO_SIGNED(-60,11),
TO_SIGNED(-13,11),
TO_SIGNED(34,11),
TO_SIGNED(81,11),
TO_SIGNED(128,11),
TO_SIGNED(174,11),
TO_SIGNED(219,11),
TO_SIGNED(264,11),
TO_SIGNED(307,11),
TO_SIGNED(349,11),
TO_SIGNED(390,11),
TO_SIGNED(430,11),
TO_SIGNED(467,11),
TO_SIGNED(503,11),
TO_SIGNED(537,11),
TO_SIGNED(569,11),
TO_SIGNED(598,11),
TO_SIGNED(625,11),
TO_SIGNED(650,11),
TO_SIGNED(672,11),
TO_SIGNED(692,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(730,11),
TO_SIGNED(718,11),
TO_SIGNED(703,11),
TO_SIGNED(685,11),
TO_SIGNED(665,11),
TO_SIGNED(642,11),
TO_SIGNED(616,11),
TO_SIGNED(588,11),
TO_SIGNED(558,11),
TO_SIGNED(526,11),
TO_SIGNED(491,11),
TO_SIGNED(455,11),
TO_SIGNED(416,11),
TO_SIGNED(376,11),
TO_SIGNED(335,11),
TO_SIGNED(292,11),
TO_SIGNED(248,11),
TO_SIGNED(204,11),
TO_SIGNED(158,11),
TO_SIGNED(112,11),
TO_SIGNED(65,11),
TO_SIGNED(18,11),
TO_SIGNED(-29,11),
TO_SIGNED(-76,11),
TO_SIGNED(-122,11),
TO_SIGNED(-168,11),
TO_SIGNED(-214,11),
TO_SIGNED(-259,11),
TO_SIGNED(-302,11),
TO_SIGNED(-345,11),
TO_SIGNED(-386,11),
TO_SIGNED(-425,11),
TO_SIGNED(-463,11),
TO_SIGNED(-499,11),
TO_SIGNED(-533,11),
TO_SIGNED(-565,11),
TO_SIGNED(-595,11),
TO_SIGNED(-622,11),
TO_SIGNED(-647,11),
TO_SIGNED(-670,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-721,11),
TO_SIGNED(-733,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-720,11),
TO_SIGNED(-705,11),
TO_SIGNED(-688,11),
TO_SIGNED(-667,11),
TO_SIGNED(-645,11),
TO_SIGNED(-619,11),
TO_SIGNED(-592,11),
TO_SIGNED(-562,11),
TO_SIGNED(-529,11),
TO_SIGNED(-495,11),
TO_SIGNED(-459,11),
TO_SIGNED(-421,11),
TO_SIGNED(-381,11),
TO_SIGNED(-340,11),
TO_SIGNED(-297,11),
TO_SIGNED(-254,11),
TO_SIGNED(-209,11),
TO_SIGNED(-163,11),
TO_SIGNED(-117,11),
TO_SIGNED(-70,11),
TO_SIGNED(-24,11),
TO_SIGNED(24,11),
TO_SIGNED(70,11),
TO_SIGNED(117,11),
TO_SIGNED(163,11),
TO_SIGNED(209,11),
TO_SIGNED(254,11),
TO_SIGNED(297,11),
TO_SIGNED(340,11),
TO_SIGNED(381,11),
TO_SIGNED(421,11),
TO_SIGNED(459,11),
TO_SIGNED(495,11),
TO_SIGNED(529,11),
TO_SIGNED(562,11),
TO_SIGNED(592,11),
TO_SIGNED(619,11),
TO_SIGNED(645,11),
TO_SIGNED(667,11),
TO_SIGNED(688,11),
TO_SIGNED(705,11),
TO_SIGNED(720,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(733,11),
TO_SIGNED(721,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(670,11),
TO_SIGNED(647,11),
TO_SIGNED(622,11),
TO_SIGNED(595,11),
TO_SIGNED(565,11),
TO_SIGNED(533,11),
TO_SIGNED(499,11),
TO_SIGNED(463,11),
TO_SIGNED(425,11),
TO_SIGNED(386,11),
TO_SIGNED(345,11),
TO_SIGNED(302,11),
TO_SIGNED(259,11),
TO_SIGNED(214,11),
TO_SIGNED(168,11),
TO_SIGNED(122,11),
TO_SIGNED(76,11),
TO_SIGNED(29,11),
TO_SIGNED(-18,11),
TO_SIGNED(-65,11),
TO_SIGNED(-112,11),
TO_SIGNED(-158,11),
TO_SIGNED(-204,11),
TO_SIGNED(-248,11),
TO_SIGNED(-292,11),
TO_SIGNED(-335,11),
TO_SIGNED(-376,11),
TO_SIGNED(-416,11),
TO_SIGNED(-455,11),
TO_SIGNED(-491,11),
TO_SIGNED(-526,11),
TO_SIGNED(-558,11),
TO_SIGNED(-588,11),
TO_SIGNED(-616,11),
TO_SIGNED(-642,11),
TO_SIGNED(-665,11),
TO_SIGNED(-685,11),
TO_SIGNED(-703,11),
TO_SIGNED(-718,11),
TO_SIGNED(-730,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-692,11),
TO_SIGNED(-672,11),
TO_SIGNED(-650,11),
TO_SIGNED(-625,11),
TO_SIGNED(-598,11),
TO_SIGNED(-569,11),
TO_SIGNED(-537,11),
TO_SIGNED(-503,11),
TO_SIGNED(-467,11),
TO_SIGNED(-430,11),
TO_SIGNED(-390,11),
TO_SIGNED(-349,11),
TO_SIGNED(-307,11),
TO_SIGNED(-264,11),
TO_SIGNED(-219,11),
TO_SIGNED(-174,11),
TO_SIGNED(-128,11),
TO_SIGNED(-81,11),
TO_SIGNED(-34,11),
TO_SIGNED(13,11),
TO_SIGNED(60,11),
TO_SIGNED(106,11),
TO_SIGNED(153,11),
TO_SIGNED(198,11),
TO_SIGNED(243,11),
TO_SIGNED(287,11),
TO_SIGNED(330,11),
TO_SIGNED(372,11),
TO_SIGNED(412,11),
TO_SIGNED(450,11),
TO_SIGNED(487,11),
TO_SIGNED(522,11),
TO_SIGNED(554,11),
TO_SIGNED(585,11),
TO_SIGNED(613,11),
TO_SIGNED(639,11),
TO_SIGNED(662,11),
TO_SIGNED(683,11),
TO_SIGNED(701,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(724,11),
TO_SIGNED(710,11),
TO_SIGNED(694,11),
TO_SIGNED(675,11),
TO_SIGNED(653,11),
TO_SIGNED(628,11),
TO_SIGNED(601,11),
TO_SIGNED(572,11),
TO_SIGNED(541,11),
TO_SIGNED(507,11),
TO_SIGNED(471,11),
TO_SIGNED(434,11),
TO_SIGNED(395,11),
TO_SIGNED(354,11),
TO_SIGNED(312,11),
TO_SIGNED(269,11),
TO_SIGNED(224,11),
TO_SIGNED(179,11),
TO_SIGNED(133,11),
TO_SIGNED(86,11),
TO_SIGNED(40,11),
TO_SIGNED(-7,11),
TO_SIGNED(-54,11),
TO_SIGNED(-101,11),
TO_SIGNED(-148,11),
TO_SIGNED(-193,11),
TO_SIGNED(-238,11),
TO_SIGNED(-282,11),
TO_SIGNED(-325,11),
TO_SIGNED(-367,11),
TO_SIGNED(-407,11),
TO_SIGNED(-446,11),
TO_SIGNED(-483,11),
TO_SIGNED(-518,11),
TO_SIGNED(-551,11),
TO_SIGNED(-582,11),
TO_SIGNED(-610,11),
TO_SIGNED(-636,11),
TO_SIGNED(-660,11),
TO_SIGNED(-681,11),
TO_SIGNED(-699,11),
TO_SIGNED(-715,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-736,11),
TO_SIGNED(-725,11),
TO_SIGNED(-712,11),
TO_SIGNED(-696,11),
TO_SIGNED(-677,11),
TO_SIGNED(-655,11),
TO_SIGNED(-631,11),
TO_SIGNED(-605,11),
TO_SIGNED(-576,11),
TO_SIGNED(-544,11),
TO_SIGNED(-511,11),
TO_SIGNED(-476,11),
TO_SIGNED(-438,11),
TO_SIGNED(-399,11),
TO_SIGNED(-359,11),
TO_SIGNED(-317,11),
TO_SIGNED(-274,11),
TO_SIGNED(-229,11),
TO_SIGNED(-184,11),
TO_SIGNED(-138,11),
TO_SIGNED(-92,11),
TO_SIGNED(-45,11),
TO_SIGNED(2,11),
TO_SIGNED(49,11),
TO_SIGNED(96,11),
TO_SIGNED(142,11),
TO_SIGNED(188,11),
TO_SIGNED(233,11),
TO_SIGNED(277,11),
TO_SIGNED(321,11),
TO_SIGNED(362,11),
TO_SIGNED(403,11),
TO_SIGNED(442,11),
TO_SIGNED(479,11),
TO_SIGNED(514,11),
TO_SIGNED(547,11),
TO_SIGNED(578,11),
TO_SIGNED(607,11),
TO_SIGNED(633,11),
TO_SIGNED(657,11),
TO_SIGNED(679,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(698,11),
TO_SIGNED(679,11),
TO_SIGNED(658,11),
TO_SIGNED(634,11),
TO_SIGNED(608,11),
TO_SIGNED(579,11),
TO_SIGNED(548,11),
TO_SIGNED(515,11),
TO_SIGNED(480,11),
TO_SIGNED(443,11),
TO_SIGNED(404,11),
TO_SIGNED(363,11),
TO_SIGNED(322,11),
TO_SIGNED(278,11),
TO_SIGNED(234,11),
TO_SIGNED(189,11),
TO_SIGNED(143,11),
TO_SIGNED(97,11),
TO_SIGNED(50,11),
TO_SIGNED(3,11),
TO_SIGNED(-44,11),
TO_SIGNED(-91,11),
TO_SIGNED(-137,11),
TO_SIGNED(-183,11),
TO_SIGNED(-228,11),
TO_SIGNED(-273,11),
TO_SIGNED(-316,11),
TO_SIGNED(-358,11),
TO_SIGNED(-398,11),
TO_SIGNED(-437,11),
TO_SIGNED(-475,11),
TO_SIGNED(-510,11),
TO_SIGNED(-544,11),
TO_SIGNED(-575,11),
TO_SIGNED(-604,11),
TO_SIGNED(-631,11),
TO_SIGNED(-655,11),
TO_SIGNED(-676,11),
TO_SIGNED(-695,11),
TO_SIGNED(-712,11),
TO_SIGNED(-725,11),
TO_SIGNED(-736,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-715,11),
TO_SIGNED(-700,11),
TO_SIGNED(-681,11),
TO_SIGNED(-660,11),
TO_SIGNED(-637,11),
TO_SIGNED(-611,11),
TO_SIGNED(-582,11),
TO_SIGNED(-552,11),
TO_SIGNED(-519,11),
TO_SIGNED(-484,11),
TO_SIGNED(-447,11),
TO_SIGNED(-408,11),
TO_SIGNED(-368,11),
TO_SIGNED(-326,11),
TO_SIGNED(-283,11),
TO_SIGNED(-239,11),
TO_SIGNED(-194,11),
TO_SIGNED(-149,11),
TO_SIGNED(-102,11),
TO_SIGNED(-56,11),
TO_SIGNED(-9,11),
TO_SIGNED(38,11),
TO_SIGNED(85,11),
TO_SIGNED(132,11),
TO_SIGNED(178,11),
TO_SIGNED(223,11),
TO_SIGNED(268,11),
TO_SIGNED(311,11),
TO_SIGNED(353,11),
TO_SIGNED(394,11),
TO_SIGNED(433,11),
TO_SIGNED(471,11),
TO_SIGNED(506,11),
TO_SIGNED(540,11),
TO_SIGNED(571,11),
TO_SIGNED(601,11),
TO_SIGNED(628,11),
TO_SIGNED(652,11),
TO_SIGNED(674,11),
TO_SIGNED(693,11),
TO_SIGNED(710,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(739,11),
TO_SIGNED(729,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(684,11),
TO_SIGNED(663,11),
TO_SIGNED(640,11),
TO_SIGNED(614,11),
TO_SIGNED(586,11),
TO_SIGNED(555,11),
TO_SIGNED(523,11),
TO_SIGNED(488,11),
TO_SIGNED(451,11),
TO_SIGNED(413,11),
TO_SIGNED(373,11),
TO_SIGNED(331,11),
TO_SIGNED(288,11),
TO_SIGNED(244,11),
TO_SIGNED(200,11),
TO_SIGNED(154,11),
TO_SIGNED(108,11),
TO_SIGNED(61,11),
TO_SIGNED(14,11),
TO_SIGNED(-33,11),
TO_SIGNED(-80,11),
TO_SIGNED(-127,11),
TO_SIGNED(-173,11),
TO_SIGNED(-218,11),
TO_SIGNED(-263,11),
TO_SIGNED(-306,11),
TO_SIGNED(-348,11),
TO_SIGNED(-389,11),
TO_SIGNED(-429,11),
TO_SIGNED(-466,11),
TO_SIGNED(-502,11),
TO_SIGNED(-536,11),
TO_SIGNED(-568,11),
TO_SIGNED(-598,11),
TO_SIGNED(-625,11),
TO_SIGNED(-650,11),
TO_SIGNED(-672,11),
TO_SIGNED(-691,11),
TO_SIGNED(-708,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-686,11),
TO_SIGNED(-665,11),
TO_SIGNED(-642,11),
TO_SIGNED(-617,11),
TO_SIGNED(-589,11),
TO_SIGNED(-559,11),
TO_SIGNED(-526,11),
TO_SIGNED(-492,11),
TO_SIGNED(-455,11),
TO_SIGNED(-417,11),
TO_SIGNED(-377,11),
TO_SIGNED(-336,11),
TO_SIGNED(-293,11),
TO_SIGNED(-249,11),
TO_SIGNED(-205,11),
TO_SIGNED(-159,11),
TO_SIGNED(-113,11),
TO_SIGNED(-66,11),
TO_SIGNED(-19,11),
TO_SIGNED(28,11),
TO_SIGNED(75,11),
TO_SIGNED(121,11),
TO_SIGNED(167,11),
TO_SIGNED(213,11),
TO_SIGNED(258,11),
TO_SIGNED(301,11),
TO_SIGNED(344,11),
TO_SIGNED(385,11),
TO_SIGNED(424,11),
TO_SIGNED(462,11),
TO_SIGNED(498,11),
TO_SIGNED(532,11),
TO_SIGNED(564,11),
TO_SIGNED(594,11),
TO_SIGNED(622,11),
TO_SIGNED(647,11),
TO_SIGNED(669,11),
TO_SIGNED(689,11),
TO_SIGNED(706,11),
TO_SIGNED(721,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(720,11),
TO_SIGNED(705,11),
TO_SIGNED(688,11),
TO_SIGNED(668,11),
TO_SIGNED(645,11),
TO_SIGNED(620,11),
TO_SIGNED(592,11),
TO_SIGNED(562,11),
TO_SIGNED(530,11),
TO_SIGNED(496,11),
TO_SIGNED(460,11),
TO_SIGNED(422,11),
TO_SIGNED(382,11),
TO_SIGNED(341,11),
TO_SIGNED(298,11),
TO_SIGNED(255,11),
TO_SIGNED(210,11),
TO_SIGNED(164,11),
TO_SIGNED(118,11),
TO_SIGNED(71,11),
TO_SIGNED(25,11),
TO_SIGNED(-22,11),
TO_SIGNED(-69,11),
TO_SIGNED(-116,11),
TO_SIGNED(-162,11),
TO_SIGNED(-208,11),
TO_SIGNED(-252,11),
TO_SIGNED(-296,11),
TO_SIGNED(-339,11),
TO_SIGNED(-380,11),
TO_SIGNED(-420,11),
TO_SIGNED(-458,11),
TO_SIGNED(-494,11),
TO_SIGNED(-529,11),
TO_SIGNED(-561,11),
TO_SIGNED(-591,11),
TO_SIGNED(-619,11),
TO_SIGNED(-644,11),
TO_SIGNED(-667,11),
TO_SIGNED(-687,11),
TO_SIGNED(-705,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-733,11),
TO_SIGNED(-721,11),
TO_SIGNED(-707,11),
TO_SIGNED(-690,11),
TO_SIGNED(-670,11),
TO_SIGNED(-648,11),
TO_SIGNED(-623,11),
TO_SIGNED(-596,11),
TO_SIGNED(-566,11),
TO_SIGNED(-534,11),
TO_SIGNED(-500,11),
TO_SIGNED(-464,11),
TO_SIGNED(-426,11),
TO_SIGNED(-387,11),
TO_SIGNED(-345,11),
TO_SIGNED(-303,11),
TO_SIGNED(-260,11),
TO_SIGNED(-215,11),
TO_SIGNED(-169,11),
TO_SIGNED(-123,11),
TO_SIGNED(-77,11),
TO_SIGNED(-30,11),
TO_SIGNED(17,11),
TO_SIGNED(64,11),
TO_SIGNED(111,11),
TO_SIGNED(157,11),
TO_SIGNED(203,11),
TO_SIGNED(247,11),
TO_SIGNED(291,11),
TO_SIGNED(334,11),
TO_SIGNED(375,11),
TO_SIGNED(415,11),
TO_SIGNED(454,11),
TO_SIGNED(490,11),
TO_SIGNED(525,11),
TO_SIGNED(557,11),
TO_SIGNED(588,11),
TO_SIGNED(616,11),
TO_SIGNED(641,11),
TO_SIGNED(664,11),
TO_SIGNED(685,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(709,11),
TO_SIGNED(692,11),
TO_SIGNED(673,11),
TO_SIGNED(651,11),
TO_SIGNED(626,11),
TO_SIGNED(599,11),
TO_SIGNED(569,11),
TO_SIGNED(538,11),
TO_SIGNED(504,11),
TO_SIGNED(468,11),
TO_SIGNED(430,11),
TO_SIGNED(391,11),
TO_SIGNED(350,11),
TO_SIGNED(308,11),
TO_SIGNED(265,11),
TO_SIGNED(220,11),
TO_SIGNED(175,11),
TO_SIGNED(129,11),
TO_SIGNED(82,11),
TO_SIGNED(35,11),
TO_SIGNED(-12,11),
TO_SIGNED(-59,11),
TO_SIGNED(-105,11),
TO_SIGNED(-152,11),
TO_SIGNED(-197,11),
TO_SIGNED(-242,11),
TO_SIGNED(-286,11),
TO_SIGNED(-329,11),
TO_SIGNED(-371,11),
TO_SIGNED(-411,11),
TO_SIGNED(-449,11),
TO_SIGNED(-486,11),
TO_SIGNED(-521,11),
TO_SIGNED(-554,11),
TO_SIGNED(-584,11),
TO_SIGNED(-613,11),
TO_SIGNED(-639,11),
TO_SIGNED(-662,11),
TO_SIGNED(-683,11),
TO_SIGNED(-701,11),
TO_SIGNED(-716,11),
TO_SIGNED(-729,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-711,11),
TO_SIGNED(-694,11),
TO_SIGNED(-675,11),
TO_SIGNED(-653,11),
TO_SIGNED(-629,11),
TO_SIGNED(-602,11),
TO_SIGNED(-573,11),
TO_SIGNED(-541,11),
TO_SIGNED(-508,11),
TO_SIGNED(-472,11),
TO_SIGNED(-435,11),
TO_SIGNED(-396,11),
TO_SIGNED(-355,11),
TO_SIGNED(-313,11),
TO_SIGNED(-270,11),
TO_SIGNED(-225,11),
TO_SIGNED(-180,11),
TO_SIGNED(-134,11),
TO_SIGNED(-87,11),
TO_SIGNED(-41,11),
TO_SIGNED(6,11),
TO_SIGNED(53,11),
TO_SIGNED(100,11),
TO_SIGNED(147,11),
TO_SIGNED(192,11),
TO_SIGNED(237,11),
TO_SIGNED(281,11),
TO_SIGNED(324,11),
TO_SIGNED(366,11),
TO_SIGNED(406,11),
TO_SIGNED(445,11),
TO_SIGNED(482,11),
TO_SIGNED(517,11),
TO_SIGNED(550,11),
TO_SIGNED(581,11),
TO_SIGNED(610,11),
TO_SIGNED(636,11),
TO_SIGNED(659,11),
TO_SIGNED(681,11),
TO_SIGNED(699,11),
TO_SIGNED(715,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(712,11),
TO_SIGNED(696,11),
TO_SIGNED(677,11),
TO_SIGNED(656,11),
TO_SIGNED(632,11),
TO_SIGNED(605,11),
TO_SIGNED(576,11),
TO_SIGNED(545,11),
TO_SIGNED(512,11),
TO_SIGNED(476,11),
TO_SIGNED(439,11),
TO_SIGNED(400,11),
TO_SIGNED(360,11),
TO_SIGNED(318,11),
TO_SIGNED(275,11),
TO_SIGNED(230,11),
TO_SIGNED(185,11),
TO_SIGNED(139,11),
TO_SIGNED(93,11),
TO_SIGNED(46,11),
TO_SIGNED(-1,11),
TO_SIGNED(-48,11),
TO_SIGNED(-95,11),
TO_SIGNED(-141,11),
TO_SIGNED(-187,11),
TO_SIGNED(-232,11),
TO_SIGNED(-276,11),
TO_SIGNED(-320,11),
TO_SIGNED(-362,11),
TO_SIGNED(-402,11),
TO_SIGNED(-441,11),
TO_SIGNED(-478,11),
TO_SIGNED(-513,11),
TO_SIGNED(-547,11),
TO_SIGNED(-578,11),
TO_SIGNED(-606,11),
TO_SIGNED(-633,11),
TO_SIGNED(-657,11),
TO_SIGNED(-678,11),
TO_SIGNED(-697,11),
TO_SIGNED(-713,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-714,11),
TO_SIGNED(-698,11),
TO_SIGNED(-680,11),
TO_SIGNED(-658,11),
TO_SIGNED(-635,11),
TO_SIGNED(-608,11),
TO_SIGNED(-580,11),
TO_SIGNED(-549,11),
TO_SIGNED(-516,11),
TO_SIGNED(-480,11),
TO_SIGNED(-443,11),
TO_SIGNED(-405,11),
TO_SIGNED(-364,11),
TO_SIGNED(-323,11),
TO_SIGNED(-279,11),
TO_SIGNED(-235,11),
TO_SIGNED(-190,11),
TO_SIGNED(-144,11),
TO_SIGNED(-98,11),
TO_SIGNED(-51,11),
TO_SIGNED(-4,11),
TO_SIGNED(43,11),
TO_SIGNED(90,11),
TO_SIGNED(136,11),
TO_SIGNED(182,11),
TO_SIGNED(227,11),
TO_SIGNED(272,11),
TO_SIGNED(315,11),
TO_SIGNED(357,11),
TO_SIGNED(397,11),
TO_SIGNED(437,11),
TO_SIGNED(474,11),
TO_SIGNED(509,11),
TO_SIGNED(543,11),
TO_SIGNED(574,11),
TO_SIGNED(603,11),
TO_SIGNED(630,11),
TO_SIGNED(654,11),
TO_SIGNED(676,11),
TO_SIGNED(695,11),
TO_SIGNED(711,11),
TO_SIGNED(725,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(716,11),
TO_SIGNED(700,11),
TO_SIGNED(682,11),
TO_SIGNED(661,11),
TO_SIGNED(637,11),
TO_SIGNED(611,11),
TO_SIGNED(583,11),
TO_SIGNED(552,11),
TO_SIGNED(519,11),
TO_SIGNED(485,11),
TO_SIGNED(448,11),
TO_SIGNED(409,11),
TO_SIGNED(369,11),
TO_SIGNED(327,11),
TO_SIGNED(284,11),
TO_SIGNED(240,11),
TO_SIGNED(195,11),
TO_SIGNED(150,11),
TO_SIGNED(103,11),
TO_SIGNED(57,11),
TO_SIGNED(10,11),
TO_SIGNED(-37,11),
TO_SIGNED(-84,11),
TO_SIGNED(-131,11),
TO_SIGNED(-177,11),
TO_SIGNED(-222,11),
TO_SIGNED(-267,11),
TO_SIGNED(-310,11),
TO_SIGNED(-352,11),
TO_SIGNED(-393,11),
TO_SIGNED(-432,11),
TO_SIGNED(-470,11),
TO_SIGNED(-505,11),
TO_SIGNED(-539,11),
TO_SIGNED(-571,11),
TO_SIGNED(-600,11),
TO_SIGNED(-627,11),
TO_SIGNED(-652,11),
TO_SIGNED(-674,11),
TO_SIGNED(-693,11),
TO_SIGNED(-710,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-702,11),
TO_SIGNED(-684,11),
TO_SIGNED(-663,11),
TO_SIGNED(-640,11),
TO_SIGNED(-615,11),
TO_SIGNED(-586,11),
TO_SIGNED(-556,11),
TO_SIGNED(-523,11),
TO_SIGNED(-489,11),
TO_SIGNED(-452,11),
TO_SIGNED(-414,11),
TO_SIGNED(-374,11),
TO_SIGNED(-332,11),
TO_SIGNED(-289,11),
TO_SIGNED(-245,11),
TO_SIGNED(-201,11),
TO_SIGNED(-155,11),
TO_SIGNED(-109,11),
TO_SIGNED(-62,11),
TO_SIGNED(-15,11),
TO_SIGNED(32,11),
TO_SIGNED(79,11),
TO_SIGNED(125,11),
TO_SIGNED(172,11),
TO_SIGNED(217,11),
TO_SIGNED(262,11),
TO_SIGNED(305,11),
TO_SIGNED(347,11),
TO_SIGNED(388,11),
TO_SIGNED(428,11),
TO_SIGNED(466,11),
TO_SIGNED(501,11),
TO_SIGNED(535,11),
TO_SIGNED(567,11),
TO_SIGNED(597,11),
TO_SIGNED(624,11),
TO_SIGNED(649,11),
TO_SIGNED(671,11),
TO_SIGNED(691,11),
TO_SIGNED(708,11),
TO_SIGNED(722,11),
TO_SIGNED(733,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(704,11),
TO_SIGNED(686,11),
TO_SIGNED(666,11),
TO_SIGNED(643,11),
TO_SIGNED(618,11),
TO_SIGNED(590,11),
TO_SIGNED(559,11),
TO_SIGNED(527,11),
TO_SIGNED(493,11),
TO_SIGNED(456,11),
TO_SIGNED(418,11),
TO_SIGNED(378,11),
TO_SIGNED(337,11),
TO_SIGNED(294,11),
TO_SIGNED(250,11),
TO_SIGNED(206,11),
TO_SIGNED(160,11),
TO_SIGNED(114,11),
TO_SIGNED(67,11),
TO_SIGNED(20,11),
TO_SIGNED(-27,11),
TO_SIGNED(-74,11),
TO_SIGNED(-120,11),
TO_SIGNED(-166,11),
TO_SIGNED(-212,11),
TO_SIGNED(-257,11),
TO_SIGNED(-300,11),
TO_SIGNED(-343,11),
TO_SIGNED(-384,11),
TO_SIGNED(-423,11),
TO_SIGNED(-461,11),
TO_SIGNED(-497,11),
TO_SIGNED(-532,11),
TO_SIGNED(-564,11),
TO_SIGNED(-594,11),
TO_SIGNED(-621,11),
TO_SIGNED(-646,11),
TO_SIGNED(-669,11),
TO_SIGNED(-689,11),
TO_SIGNED(-706,11),
TO_SIGNED(-721,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-720,11),
TO_SIGNED(-706,11),
TO_SIGNED(-688,11),
TO_SIGNED(-668,11),
TO_SIGNED(-646,11),
TO_SIGNED(-621,11),
TO_SIGNED(-593,11),
TO_SIGNED(-563,11),
TO_SIGNED(-531,11),
TO_SIGNED(-497,11),
TO_SIGNED(-460,11),
TO_SIGNED(-422,11),
TO_SIGNED(-383,11),
TO_SIGNED(-342,11),
TO_SIGNED(-299,11),
TO_SIGNED(-256,11),
TO_SIGNED(-211,11),
TO_SIGNED(-165,11),
TO_SIGNED(-119,11),
TO_SIGNED(-73,11),
TO_SIGNED(-26,11),
TO_SIGNED(21,11),
TO_SIGNED(68,11),
TO_SIGNED(115,11),
TO_SIGNED(161,11),
TO_SIGNED(207,11),
TO_SIGNED(251,11),
TO_SIGNED(295,11),
TO_SIGNED(338,11),
TO_SIGNED(379,11),
TO_SIGNED(419,11),
TO_SIGNED(457,11),
TO_SIGNED(493,11),
TO_SIGNED(528,11),
TO_SIGNED(560,11),
TO_SIGNED(590,11),
TO_SIGNED(618,11),
TO_SIGNED(644,11),
TO_SIGNED(666,11),
TO_SIGNED(687,11),
TO_SIGNED(704,11),
TO_SIGNED(719,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(671,11),
TO_SIGNED(648,11),
TO_SIGNED(624,11),
TO_SIGNED(596,11),
TO_SIGNED(567,11),
TO_SIGNED(535,11),
TO_SIGNED(501,11),
TO_SIGNED(465,11),
TO_SIGNED(427,11),
TO_SIGNED(387,11),
TO_SIGNED(346,11),
TO_SIGNED(304,11),
TO_SIGNED(261,11),
TO_SIGNED(216,11),
TO_SIGNED(171,11),
TO_SIGNED(124,11),
TO_SIGNED(78,11),
TO_SIGNED(31,11),
TO_SIGNED(-16,11),
TO_SIGNED(-63,11),
TO_SIGNED(-110,11),
TO_SIGNED(-156,11),
TO_SIGNED(-202,11),
TO_SIGNED(-246,11),
TO_SIGNED(-290,11),
TO_SIGNED(-333,11),
TO_SIGNED(-375,11),
TO_SIGNED(-415,11),
TO_SIGNED(-453,11),
TO_SIGNED(-489,11),
TO_SIGNED(-524,11),
TO_SIGNED(-557,11),
TO_SIGNED(-587,11),
TO_SIGNED(-615,11),
TO_SIGNED(-641,11),
TO_SIGNED(-664,11),
TO_SIGNED(-685,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-730,11),
TO_SIGNED(-739,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-693,11),
TO_SIGNED(-673,11),
TO_SIGNED(-651,11),
TO_SIGNED(-627,11),
TO_SIGNED(-599,11),
TO_SIGNED(-570,11),
TO_SIGNED(-538,11),
TO_SIGNED(-505,11),
TO_SIGNED(-469,11),
TO_SIGNED(-431,11),
TO_SIGNED(-392,11),
TO_SIGNED(-351,11),
TO_SIGNED(-309,11),
TO_SIGNED(-266,11),
TO_SIGNED(-221,11),
TO_SIGNED(-176,11),
TO_SIGNED(-130,11),
TO_SIGNED(-83,11),
TO_SIGNED(-36,11),
TO_SIGNED(11,11),
TO_SIGNED(58,11),
TO_SIGNED(104,11),
TO_SIGNED(151,11),
TO_SIGNED(196,11),
TO_SIGNED(241,11),
TO_SIGNED(285,11),
TO_SIGNED(328,11),
TO_SIGNED(370,11),
TO_SIGNED(410,11),
TO_SIGNED(449,11),
TO_SIGNED(485,11),
TO_SIGNED(520,11),
TO_SIGNED(553,11),
TO_SIGNED(584,11),
TO_SIGNED(612,11),
TO_SIGNED(638,11),
TO_SIGNED(661,11),
TO_SIGNED(682,11),
TO_SIGNED(700,11),
TO_SIGNED(716,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(725,11),
TO_SIGNED(711,11),
TO_SIGNED(695,11),
TO_SIGNED(675,11),
TO_SIGNED(654,11),
TO_SIGNED(629,11),
TO_SIGNED(603,11),
TO_SIGNED(574,11),
TO_SIGNED(542,11),
TO_SIGNED(509,11),
TO_SIGNED(473,11),
TO_SIGNED(436,11),
TO_SIGNED(397,11),
TO_SIGNED(356,11),
TO_SIGNED(314,11),
TO_SIGNED(271,11),
TO_SIGNED(226,11),
TO_SIGNED(181,11),
TO_SIGNED(135,11),
TO_SIGNED(88,11),
TO_SIGNED(42,11),
TO_SIGNED(-5,11),
TO_SIGNED(-52,11),
TO_SIGNED(-99,11),
TO_SIGNED(-145,11),
TO_SIGNED(-191,11),
TO_SIGNED(-236,11),
TO_SIGNED(-280,11),
TO_SIGNED(-323,11),
TO_SIGNED(-365,11),
TO_SIGNED(-406,11),
TO_SIGNED(-444,11),
TO_SIGNED(-481,11),
TO_SIGNED(-516,11),
TO_SIGNED(-549,11),
TO_SIGNED(-580,11),
TO_SIGNED(-609,11),
TO_SIGNED(-635,11),
TO_SIGNED(-659,11),
TO_SIGNED(-680,11),
TO_SIGNED(-699,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-736,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-678,11),
TO_SIGNED(-656,11),
TO_SIGNED(-632,11),
TO_SIGNED(-606,11),
TO_SIGNED(-577,11),
TO_SIGNED(-546,11),
TO_SIGNED(-512,11),
TO_SIGNED(-477,11),
TO_SIGNED(-440,11),
TO_SIGNED(-401,11),
TO_SIGNED(-361,11),
TO_SIGNED(-319,11),
TO_SIGNED(-275,11),
TO_SIGNED(-231,11),
TO_SIGNED(-186,11),
TO_SIGNED(-140,11),
TO_SIGNED(-94,11),
TO_SIGNED(-47,11),
TO_SIGNED(0,11),
TO_SIGNED(47,11),
TO_SIGNED(94,11),
TO_SIGNED(140,11),
TO_SIGNED(186,11),
TO_SIGNED(231,11),
TO_SIGNED(275,11),
TO_SIGNED(319,11),
TO_SIGNED(361,11),
TO_SIGNED(401,11),
TO_SIGNED(440,11),
TO_SIGNED(477,11),
TO_SIGNED(512,11),
TO_SIGNED(546,11),
TO_SIGNED(577,11),
TO_SIGNED(606,11),
TO_SIGNED(632,11),
TO_SIGNED(656,11),
TO_SIGNED(678,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(736,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(699,11),
TO_SIGNED(680,11),
TO_SIGNED(659,11),
TO_SIGNED(635,11),
TO_SIGNED(609,11),
TO_SIGNED(580,11),
TO_SIGNED(549,11),
TO_SIGNED(516,11),
TO_SIGNED(481,11),
TO_SIGNED(444,11),
TO_SIGNED(406,11),
TO_SIGNED(365,11),
TO_SIGNED(323,11),
TO_SIGNED(280,11),
TO_SIGNED(236,11),
TO_SIGNED(191,11),
TO_SIGNED(145,11),
TO_SIGNED(99,11),
TO_SIGNED(52,11),
TO_SIGNED(5,11),
TO_SIGNED(-42,11),
TO_SIGNED(-88,11),
TO_SIGNED(-135,11),
TO_SIGNED(-181,11),
TO_SIGNED(-226,11),
TO_SIGNED(-271,11),
TO_SIGNED(-314,11),
TO_SIGNED(-356,11),
TO_SIGNED(-397,11),
TO_SIGNED(-436,11),
TO_SIGNED(-473,11),
TO_SIGNED(-509,11),
TO_SIGNED(-542,11),
TO_SIGNED(-574,11),
TO_SIGNED(-603,11),
TO_SIGNED(-629,11),
TO_SIGNED(-654,11),
TO_SIGNED(-675,11),
TO_SIGNED(-695,11),
TO_SIGNED(-711,11),
TO_SIGNED(-725,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-716,11),
TO_SIGNED(-700,11),
TO_SIGNED(-682,11),
TO_SIGNED(-661,11),
TO_SIGNED(-638,11),
TO_SIGNED(-612,11),
TO_SIGNED(-584,11),
TO_SIGNED(-553,11),
TO_SIGNED(-520,11),
TO_SIGNED(-485,11),
TO_SIGNED(-449,11),
TO_SIGNED(-410,11),
TO_SIGNED(-370,11),
TO_SIGNED(-328,11),
TO_SIGNED(-285,11),
TO_SIGNED(-241,11),
TO_SIGNED(-196,11),
TO_SIGNED(-151,11),
TO_SIGNED(-104,11),
TO_SIGNED(-58,11),
TO_SIGNED(-11,11),
TO_SIGNED(36,11),
TO_SIGNED(83,11),
TO_SIGNED(130,11),
TO_SIGNED(176,11),
TO_SIGNED(221,11),
TO_SIGNED(266,11),
TO_SIGNED(309,11),
TO_SIGNED(351,11),
TO_SIGNED(392,11),
TO_SIGNED(431,11),
TO_SIGNED(469,11),
TO_SIGNED(505,11),
TO_SIGNED(538,11),
TO_SIGNED(570,11),
TO_SIGNED(599,11),
TO_SIGNED(627,11),
TO_SIGNED(651,11),
TO_SIGNED(673,11),
TO_SIGNED(693,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(739,11),
TO_SIGNED(730,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(685,11),
TO_SIGNED(664,11),
TO_SIGNED(641,11),
TO_SIGNED(615,11),
TO_SIGNED(587,11),
TO_SIGNED(557,11),
TO_SIGNED(524,11),
TO_SIGNED(489,11),
TO_SIGNED(453,11),
TO_SIGNED(415,11),
TO_SIGNED(375,11),
TO_SIGNED(333,11),
TO_SIGNED(290,11),
TO_SIGNED(246,11),
TO_SIGNED(202,11),
TO_SIGNED(156,11),
TO_SIGNED(110,11),
TO_SIGNED(63,11),
TO_SIGNED(16,11),
TO_SIGNED(-31,11),
TO_SIGNED(-78,11),
TO_SIGNED(-124,11),
TO_SIGNED(-171,11),
TO_SIGNED(-216,11),
TO_SIGNED(-261,11),
TO_SIGNED(-304,11),
TO_SIGNED(-346,11),
TO_SIGNED(-387,11),
TO_SIGNED(-427,11),
TO_SIGNED(-465,11),
TO_SIGNED(-501,11),
TO_SIGNED(-535,11),
TO_SIGNED(-567,11),
TO_SIGNED(-596,11),
TO_SIGNED(-624,11),
TO_SIGNED(-648,11),
TO_SIGNED(-671,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-719,11),
TO_SIGNED(-704,11),
TO_SIGNED(-687,11),
TO_SIGNED(-666,11),
TO_SIGNED(-644,11),
TO_SIGNED(-618,11),
TO_SIGNED(-590,11),
TO_SIGNED(-560,11),
TO_SIGNED(-528,11),
TO_SIGNED(-493,11),
TO_SIGNED(-457,11),
TO_SIGNED(-419,11),
TO_SIGNED(-379,11),
TO_SIGNED(-338,11),
TO_SIGNED(-295,11),
TO_SIGNED(-251,11),
TO_SIGNED(-207,11),
TO_SIGNED(-161,11),
TO_SIGNED(-115,11),
TO_SIGNED(-68,11),
TO_SIGNED(-21,11),
TO_SIGNED(26,11),
TO_SIGNED(73,11),
TO_SIGNED(119,11),
TO_SIGNED(165,11),
TO_SIGNED(211,11),
TO_SIGNED(256,11),
TO_SIGNED(299,11),
TO_SIGNED(342,11),
TO_SIGNED(383,11),
TO_SIGNED(422,11),
TO_SIGNED(460,11),
TO_SIGNED(497,11),
TO_SIGNED(531,11),
TO_SIGNED(563,11),
TO_SIGNED(593,11),
TO_SIGNED(621,11),
TO_SIGNED(646,11),
TO_SIGNED(668,11),
TO_SIGNED(688,11),
TO_SIGNED(706,11),
TO_SIGNED(720,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(721,11),
TO_SIGNED(706,11),
TO_SIGNED(689,11),
TO_SIGNED(669,11),
TO_SIGNED(646,11),
TO_SIGNED(621,11),
TO_SIGNED(594,11),
TO_SIGNED(564,11),
TO_SIGNED(532,11),
TO_SIGNED(497,11),
TO_SIGNED(461,11),
TO_SIGNED(423,11),
TO_SIGNED(384,11),
TO_SIGNED(343,11),
TO_SIGNED(300,11),
TO_SIGNED(257,11),
TO_SIGNED(212,11),
TO_SIGNED(166,11),
TO_SIGNED(120,11),
TO_SIGNED(74,11),
TO_SIGNED(27,11),
TO_SIGNED(-20,11),
TO_SIGNED(-67,11),
TO_SIGNED(-114,11),
TO_SIGNED(-160,11),
TO_SIGNED(-206,11),
TO_SIGNED(-250,11),
TO_SIGNED(-294,11),
TO_SIGNED(-337,11),
TO_SIGNED(-378,11),
TO_SIGNED(-418,11),
TO_SIGNED(-456,11),
TO_SIGNED(-493,11),
TO_SIGNED(-527,11),
TO_SIGNED(-559,11),
TO_SIGNED(-590,11),
TO_SIGNED(-618,11),
TO_SIGNED(-643,11),
TO_SIGNED(-666,11),
TO_SIGNED(-686,11),
TO_SIGNED(-704,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-733,11),
TO_SIGNED(-722,11),
TO_SIGNED(-708,11),
TO_SIGNED(-691,11),
TO_SIGNED(-671,11),
TO_SIGNED(-649,11),
TO_SIGNED(-624,11),
TO_SIGNED(-597,11),
TO_SIGNED(-567,11),
TO_SIGNED(-535,11),
TO_SIGNED(-501,11),
TO_SIGNED(-466,11),
TO_SIGNED(-428,11),
TO_SIGNED(-388,11),
TO_SIGNED(-347,11),
TO_SIGNED(-305,11),
TO_SIGNED(-262,11),
TO_SIGNED(-217,11),
TO_SIGNED(-172,11),
TO_SIGNED(-125,11),
TO_SIGNED(-79,11),
TO_SIGNED(-32,11),
TO_SIGNED(15,11),
TO_SIGNED(62,11),
TO_SIGNED(109,11),
TO_SIGNED(155,11),
TO_SIGNED(201,11),
TO_SIGNED(245,11),
TO_SIGNED(289,11),
TO_SIGNED(332,11),
TO_SIGNED(374,11),
TO_SIGNED(414,11),
TO_SIGNED(452,11),
TO_SIGNED(489,11),
TO_SIGNED(523,11),
TO_SIGNED(556,11),
TO_SIGNED(586,11),
TO_SIGNED(615,11),
TO_SIGNED(640,11),
TO_SIGNED(663,11),
TO_SIGNED(684,11),
TO_SIGNED(702,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(710,11),
TO_SIGNED(693,11),
TO_SIGNED(674,11),
TO_SIGNED(652,11),
TO_SIGNED(627,11),
TO_SIGNED(600,11),
TO_SIGNED(571,11),
TO_SIGNED(539,11),
TO_SIGNED(505,11),
TO_SIGNED(470,11),
TO_SIGNED(432,11),
TO_SIGNED(393,11),
TO_SIGNED(352,11),
TO_SIGNED(310,11),
TO_SIGNED(267,11),
TO_SIGNED(222,11),
TO_SIGNED(177,11),
TO_SIGNED(131,11),
TO_SIGNED(84,11),
TO_SIGNED(37,11),
TO_SIGNED(-10,11),
TO_SIGNED(-57,11),
TO_SIGNED(-103,11),
TO_SIGNED(-150,11),
TO_SIGNED(-195,11),
TO_SIGNED(-240,11),
TO_SIGNED(-284,11),
TO_SIGNED(-327,11),
TO_SIGNED(-369,11),
TO_SIGNED(-409,11),
TO_SIGNED(-448,11),
TO_SIGNED(-485,11),
TO_SIGNED(-519,11),
TO_SIGNED(-552,11),
TO_SIGNED(-583,11),
TO_SIGNED(-611,11),
TO_SIGNED(-637,11),
TO_SIGNED(-661,11),
TO_SIGNED(-682,11),
TO_SIGNED(-700,11),
TO_SIGNED(-716,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-725,11),
TO_SIGNED(-711,11),
TO_SIGNED(-695,11),
TO_SIGNED(-676,11),
TO_SIGNED(-654,11),
TO_SIGNED(-630,11),
TO_SIGNED(-603,11),
TO_SIGNED(-574,11),
TO_SIGNED(-543,11),
TO_SIGNED(-509,11),
TO_SIGNED(-474,11),
TO_SIGNED(-437,11),
TO_SIGNED(-397,11),
TO_SIGNED(-357,11),
TO_SIGNED(-315,11),
TO_SIGNED(-272,11),
TO_SIGNED(-227,11),
TO_SIGNED(-182,11),
TO_SIGNED(-136,11),
TO_SIGNED(-90,11),
TO_SIGNED(-43,11),
TO_SIGNED(4,11),
TO_SIGNED(51,11),
TO_SIGNED(98,11),
TO_SIGNED(144,11),
TO_SIGNED(190,11),
TO_SIGNED(235,11),
TO_SIGNED(279,11),
TO_SIGNED(323,11),
TO_SIGNED(364,11),
TO_SIGNED(405,11),
TO_SIGNED(443,11),
TO_SIGNED(480,11),
TO_SIGNED(516,11),
TO_SIGNED(549,11),
TO_SIGNED(580,11),
TO_SIGNED(608,11),
TO_SIGNED(635,11),
TO_SIGNED(658,11),
TO_SIGNED(680,11),
TO_SIGNED(698,11),
TO_SIGNED(714,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(713,11),
TO_SIGNED(697,11),
TO_SIGNED(678,11),
TO_SIGNED(657,11),
TO_SIGNED(633,11),
TO_SIGNED(606,11),
TO_SIGNED(578,11),
TO_SIGNED(547,11),
TO_SIGNED(513,11),
TO_SIGNED(478,11),
TO_SIGNED(441,11),
TO_SIGNED(402,11),
TO_SIGNED(362,11),
TO_SIGNED(320,11),
TO_SIGNED(276,11),
TO_SIGNED(232,11),
TO_SIGNED(187,11),
TO_SIGNED(141,11),
TO_SIGNED(95,11),
TO_SIGNED(48,11),
TO_SIGNED(1,11),
TO_SIGNED(-46,11),
TO_SIGNED(-93,11),
TO_SIGNED(-139,11),
TO_SIGNED(-185,11),
TO_SIGNED(-230,11),
TO_SIGNED(-275,11),
TO_SIGNED(-318,11),
TO_SIGNED(-360,11),
TO_SIGNED(-400,11),
TO_SIGNED(-439,11),
TO_SIGNED(-476,11),
TO_SIGNED(-512,11),
TO_SIGNED(-545,11),
TO_SIGNED(-576,11),
TO_SIGNED(-605,11),
TO_SIGNED(-632,11),
TO_SIGNED(-656,11),
TO_SIGNED(-677,11),
TO_SIGNED(-696,11),
TO_SIGNED(-712,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-715,11),
TO_SIGNED(-699,11),
TO_SIGNED(-681,11),
TO_SIGNED(-659,11),
TO_SIGNED(-636,11),
TO_SIGNED(-610,11),
TO_SIGNED(-581,11),
TO_SIGNED(-550,11),
TO_SIGNED(-517,11),
TO_SIGNED(-482,11),
TO_SIGNED(-445,11),
TO_SIGNED(-406,11),
TO_SIGNED(-366,11),
TO_SIGNED(-324,11),
TO_SIGNED(-281,11),
TO_SIGNED(-237,11),
TO_SIGNED(-192,11),
TO_SIGNED(-147,11),
TO_SIGNED(-100,11),
TO_SIGNED(-53,11),
TO_SIGNED(-6,11),
TO_SIGNED(41,11),
TO_SIGNED(87,11),
TO_SIGNED(134,11),
TO_SIGNED(180,11),
TO_SIGNED(225,11),
TO_SIGNED(270,11),
TO_SIGNED(313,11),
TO_SIGNED(355,11),
TO_SIGNED(396,11),
TO_SIGNED(435,11),
TO_SIGNED(472,11),
TO_SIGNED(508,11),
TO_SIGNED(541,11),
TO_SIGNED(573,11),
TO_SIGNED(602,11),
TO_SIGNED(629,11),
TO_SIGNED(653,11),
TO_SIGNED(675,11),
TO_SIGNED(694,11),
TO_SIGNED(711,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(729,11),
TO_SIGNED(716,11),
TO_SIGNED(701,11),
TO_SIGNED(683,11),
TO_SIGNED(662,11),
TO_SIGNED(639,11),
TO_SIGNED(613,11),
TO_SIGNED(584,11),
TO_SIGNED(554,11),
TO_SIGNED(521,11),
TO_SIGNED(486,11),
TO_SIGNED(449,11),
TO_SIGNED(411,11),
TO_SIGNED(371,11),
TO_SIGNED(329,11),
TO_SIGNED(286,11),
TO_SIGNED(242,11),
TO_SIGNED(197,11),
TO_SIGNED(152,11),
TO_SIGNED(105,11),
TO_SIGNED(59,11),
TO_SIGNED(12,11),
TO_SIGNED(-35,11),
TO_SIGNED(-82,11),
TO_SIGNED(-129,11),
TO_SIGNED(-175,11),
TO_SIGNED(-220,11),
TO_SIGNED(-265,11),
TO_SIGNED(-308,11),
TO_SIGNED(-350,11),
TO_SIGNED(-391,11),
TO_SIGNED(-430,11),
TO_SIGNED(-468,11),
TO_SIGNED(-504,11),
TO_SIGNED(-538,11),
TO_SIGNED(-569,11),
TO_SIGNED(-599,11),
TO_SIGNED(-626,11),
TO_SIGNED(-651,11),
TO_SIGNED(-673,11),
TO_SIGNED(-692,11),
TO_SIGNED(-709,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-685,11),
TO_SIGNED(-664,11),
TO_SIGNED(-641,11),
TO_SIGNED(-616,11),
TO_SIGNED(-588,11),
TO_SIGNED(-557,11),
TO_SIGNED(-525,11),
TO_SIGNED(-490,11),
TO_SIGNED(-454,11),
TO_SIGNED(-415,11),
TO_SIGNED(-375,11),
TO_SIGNED(-334,11),
TO_SIGNED(-291,11),
TO_SIGNED(-247,11),
TO_SIGNED(-203,11),
TO_SIGNED(-157,11),
TO_SIGNED(-111,11),
TO_SIGNED(-64,11),
TO_SIGNED(-17,11),
TO_SIGNED(30,11),
TO_SIGNED(77,11),
TO_SIGNED(123,11),
TO_SIGNED(169,11),
TO_SIGNED(215,11),
TO_SIGNED(260,11),
TO_SIGNED(303,11),
TO_SIGNED(345,11),
TO_SIGNED(387,11),
TO_SIGNED(426,11),
TO_SIGNED(464,11),
TO_SIGNED(500,11),
TO_SIGNED(534,11),
TO_SIGNED(566,11),
TO_SIGNED(596,11),
TO_SIGNED(623,11),
TO_SIGNED(648,11),
TO_SIGNED(670,11),
TO_SIGNED(690,11),
TO_SIGNED(707,11),
TO_SIGNED(721,11),
TO_SIGNED(733,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(705,11),
TO_SIGNED(687,11),
TO_SIGNED(667,11),
TO_SIGNED(644,11),
TO_SIGNED(619,11),
TO_SIGNED(591,11),
TO_SIGNED(561,11),
TO_SIGNED(529,11),
TO_SIGNED(494,11),
TO_SIGNED(458,11),
TO_SIGNED(420,11),
TO_SIGNED(380,11),
TO_SIGNED(339,11),
TO_SIGNED(296,11),
TO_SIGNED(252,11),
TO_SIGNED(208,11),
TO_SIGNED(162,11),
TO_SIGNED(116,11),
TO_SIGNED(69,11),
TO_SIGNED(22,11),
TO_SIGNED(-25,11),
TO_SIGNED(-71,11),
TO_SIGNED(-118,11),
TO_SIGNED(-164,11),
TO_SIGNED(-210,11),
TO_SIGNED(-255,11),
TO_SIGNED(-298,11),
TO_SIGNED(-341,11),
TO_SIGNED(-382,11),
TO_SIGNED(-422,11),
TO_SIGNED(-460,11),
TO_SIGNED(-496,11),
TO_SIGNED(-530,11),
TO_SIGNED(-562,11),
TO_SIGNED(-592,11),
TO_SIGNED(-620,11),
TO_SIGNED(-645,11),
TO_SIGNED(-668,11),
TO_SIGNED(-688,11),
TO_SIGNED(-705,11),
TO_SIGNED(-720,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-721,11),
TO_SIGNED(-706,11),
TO_SIGNED(-689,11),
TO_SIGNED(-669,11),
TO_SIGNED(-647,11),
TO_SIGNED(-622,11),
TO_SIGNED(-594,11),
TO_SIGNED(-564,11),
TO_SIGNED(-532,11),
TO_SIGNED(-498,11),
TO_SIGNED(-462,11),
TO_SIGNED(-424,11),
TO_SIGNED(-385,11),
TO_SIGNED(-344,11),
TO_SIGNED(-301,11),
TO_SIGNED(-258,11),
TO_SIGNED(-213,11),
TO_SIGNED(-167,11),
TO_SIGNED(-121,11),
TO_SIGNED(-75,11),
TO_SIGNED(-28,11),
TO_SIGNED(19,11),
TO_SIGNED(66,11),
TO_SIGNED(113,11),
TO_SIGNED(159,11),
TO_SIGNED(205,11),
TO_SIGNED(249,11),
TO_SIGNED(293,11),
TO_SIGNED(336,11),
TO_SIGNED(377,11),
TO_SIGNED(417,11),
TO_SIGNED(455,11),
TO_SIGNED(492,11),
TO_SIGNED(526,11),
TO_SIGNED(559,11),
TO_SIGNED(589,11),
TO_SIGNED(617,11),
TO_SIGNED(642,11),
TO_SIGNED(665,11),
TO_SIGNED(686,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(708,11),
TO_SIGNED(691,11),
TO_SIGNED(672,11),
TO_SIGNED(650,11),
TO_SIGNED(625,11),
TO_SIGNED(598,11),
TO_SIGNED(568,11),
TO_SIGNED(536,11),
TO_SIGNED(502,11),
TO_SIGNED(466,11),
TO_SIGNED(429,11),
TO_SIGNED(389,11),
TO_SIGNED(348,11),
TO_SIGNED(306,11),
TO_SIGNED(263,11),
TO_SIGNED(218,11),
TO_SIGNED(173,11),
TO_SIGNED(127,11),
TO_SIGNED(80,11),
TO_SIGNED(33,11),
TO_SIGNED(-14,11),
TO_SIGNED(-61,11),
TO_SIGNED(-108,11),
TO_SIGNED(-154,11),
TO_SIGNED(-200,11),
TO_SIGNED(-244,11),
TO_SIGNED(-288,11),
TO_SIGNED(-331,11),
TO_SIGNED(-373,11),
TO_SIGNED(-413,11),
TO_SIGNED(-451,11),
TO_SIGNED(-488,11),
TO_SIGNED(-523,11),
TO_SIGNED(-555,11),
TO_SIGNED(-586,11),
TO_SIGNED(-614,11),
TO_SIGNED(-640,11),
TO_SIGNED(-663,11),
TO_SIGNED(-684,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-729,11),
TO_SIGNED(-739,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-710,11),
TO_SIGNED(-693,11),
TO_SIGNED(-674,11),
TO_SIGNED(-652,11),
TO_SIGNED(-628,11),
TO_SIGNED(-601,11),
TO_SIGNED(-571,11),
TO_SIGNED(-540,11),
TO_SIGNED(-506,11),
TO_SIGNED(-471,11),
TO_SIGNED(-433,11),
TO_SIGNED(-394,11),
TO_SIGNED(-353,11),
TO_SIGNED(-311,11),
TO_SIGNED(-268,11),
TO_SIGNED(-223,11),
TO_SIGNED(-178,11),
TO_SIGNED(-132,11),
TO_SIGNED(-85,11),
TO_SIGNED(-38,11),
TO_SIGNED(9,11),
TO_SIGNED(56,11),
TO_SIGNED(102,11),
TO_SIGNED(149,11),
TO_SIGNED(194,11),
TO_SIGNED(239,11),
TO_SIGNED(283,11),
TO_SIGNED(326,11),
TO_SIGNED(368,11),
TO_SIGNED(408,11),
TO_SIGNED(447,11),
TO_SIGNED(484,11),
TO_SIGNED(519,11),
TO_SIGNED(552,11),
TO_SIGNED(582,11),
TO_SIGNED(611,11),
TO_SIGNED(637,11),
TO_SIGNED(660,11),
TO_SIGNED(681,11),
TO_SIGNED(700,11),
TO_SIGNED(715,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(736,11),
TO_SIGNED(725,11),
TO_SIGNED(712,11),
TO_SIGNED(695,11),
TO_SIGNED(676,11),
TO_SIGNED(655,11),
TO_SIGNED(631,11),
TO_SIGNED(604,11),
TO_SIGNED(575,11),
TO_SIGNED(544,11),
TO_SIGNED(510,11),
TO_SIGNED(475,11),
TO_SIGNED(437,11),
TO_SIGNED(398,11),
TO_SIGNED(358,11),
TO_SIGNED(316,11),
TO_SIGNED(273,11),
TO_SIGNED(228,11),
TO_SIGNED(183,11),
TO_SIGNED(137,11),
TO_SIGNED(91,11),
TO_SIGNED(44,11),
TO_SIGNED(-3,11),
TO_SIGNED(-50,11),
TO_SIGNED(-97,11),
TO_SIGNED(-143,11),
TO_SIGNED(-189,11),
TO_SIGNED(-234,11),
TO_SIGNED(-278,11),
TO_SIGNED(-322,11),
TO_SIGNED(-363,11),
TO_SIGNED(-404,11),
TO_SIGNED(-443,11),
TO_SIGNED(-480,11),
TO_SIGNED(-515,11),
TO_SIGNED(-548,11),
TO_SIGNED(-579,11),
TO_SIGNED(-608,11),
TO_SIGNED(-634,11),
TO_SIGNED(-658,11),
TO_SIGNED(-679,11),
TO_SIGNED(-698,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-679,11),
TO_SIGNED(-657,11),
TO_SIGNED(-633,11),
TO_SIGNED(-607,11),
TO_SIGNED(-578,11),
TO_SIGNED(-547,11),
TO_SIGNED(-514,11),
TO_SIGNED(-479,11),
TO_SIGNED(-442,11),
TO_SIGNED(-403,11),
TO_SIGNED(-362,11),
TO_SIGNED(-321,11),
TO_SIGNED(-277,11),
TO_SIGNED(-233,11),
TO_SIGNED(-188,11),
TO_SIGNED(-142,11),
TO_SIGNED(-96,11),
TO_SIGNED(-49,11),
TO_SIGNED(-2,11),
TO_SIGNED(45,11),
TO_SIGNED(92,11),
TO_SIGNED(138,11),
TO_SIGNED(184,11),
TO_SIGNED(229,11),
TO_SIGNED(274,11),
TO_SIGNED(317,11),
TO_SIGNED(359,11),
TO_SIGNED(399,11),
TO_SIGNED(438,11),
TO_SIGNED(476,11),
TO_SIGNED(511,11),
TO_SIGNED(544,11),
TO_SIGNED(576,11),
TO_SIGNED(605,11),
TO_SIGNED(631,11),
TO_SIGNED(655,11),
TO_SIGNED(677,11),
TO_SIGNED(696,11),
TO_SIGNED(712,11),
TO_SIGNED(725,11),
TO_SIGNED(736,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(715,11),
TO_SIGNED(699,11),
TO_SIGNED(681,11),
TO_SIGNED(660,11),
TO_SIGNED(636,11),
TO_SIGNED(610,11),
TO_SIGNED(582,11),
TO_SIGNED(551,11),
TO_SIGNED(518,11),
TO_SIGNED(483,11),
TO_SIGNED(446,11),
TO_SIGNED(407,11),
TO_SIGNED(367,11),
TO_SIGNED(325,11),
TO_SIGNED(282,11),
TO_SIGNED(238,11),
TO_SIGNED(193,11),
TO_SIGNED(148,11),
TO_SIGNED(101,11),
TO_SIGNED(54,11),
TO_SIGNED(7,11),
TO_SIGNED(-40,11),
TO_SIGNED(-86,11),
TO_SIGNED(-133,11),
TO_SIGNED(-179,11),
TO_SIGNED(-224,11),
TO_SIGNED(-269,11),
TO_SIGNED(-312,11),
TO_SIGNED(-354,11),
TO_SIGNED(-395,11),
TO_SIGNED(-434,11),
TO_SIGNED(-471,11),
TO_SIGNED(-507,11),
TO_SIGNED(-541,11),
TO_SIGNED(-572,11),
TO_SIGNED(-601,11),
TO_SIGNED(-628,11),
TO_SIGNED(-653,11),
TO_SIGNED(-675,11),
TO_SIGNED(-694,11),
TO_SIGNED(-710,11),
TO_SIGNED(-724,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-701,11),
TO_SIGNED(-683,11),
TO_SIGNED(-662,11),
TO_SIGNED(-639,11),
TO_SIGNED(-613,11),
TO_SIGNED(-585,11),
TO_SIGNED(-554,11),
TO_SIGNED(-522,11),
TO_SIGNED(-487,11),
TO_SIGNED(-450,11),
TO_SIGNED(-412,11),
TO_SIGNED(-372,11),
TO_SIGNED(-330,11),
TO_SIGNED(-287,11),
TO_SIGNED(-243,11),
TO_SIGNED(-198,11),
TO_SIGNED(-153,11),
TO_SIGNED(-106,11),
TO_SIGNED(-60,11),
TO_SIGNED(-13,11),
TO_SIGNED(34,11),
TO_SIGNED(81,11),
TO_SIGNED(128,11),
TO_SIGNED(174,11),
TO_SIGNED(219,11),
TO_SIGNED(264,11),
TO_SIGNED(307,11),
TO_SIGNED(349,11),
TO_SIGNED(390,11),
TO_SIGNED(430,11),
TO_SIGNED(467,11),
TO_SIGNED(503,11),
TO_SIGNED(537,11),
TO_SIGNED(569,11),
TO_SIGNED(598,11),
TO_SIGNED(625,11),
TO_SIGNED(650,11),
TO_SIGNED(672,11),
TO_SIGNED(692,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(730,11),
TO_SIGNED(718,11),
TO_SIGNED(703,11),
TO_SIGNED(685,11),
TO_SIGNED(665,11),
TO_SIGNED(642,11),
TO_SIGNED(616,11),
TO_SIGNED(588,11),
TO_SIGNED(558,11),
TO_SIGNED(526,11),
TO_SIGNED(491,11),
TO_SIGNED(455,11),
TO_SIGNED(416,11),
TO_SIGNED(376,11),
TO_SIGNED(335,11),
TO_SIGNED(292,11),
TO_SIGNED(248,11),
TO_SIGNED(204,11),
TO_SIGNED(158,11),
TO_SIGNED(112,11),
TO_SIGNED(65,11),
TO_SIGNED(18,11),
TO_SIGNED(-29,11),
TO_SIGNED(-76,11),
TO_SIGNED(-122,11),
TO_SIGNED(-168,11),
TO_SIGNED(-214,11),
TO_SIGNED(-259,11),
TO_SIGNED(-302,11),
TO_SIGNED(-345,11),
TO_SIGNED(-386,11),
TO_SIGNED(-425,11),
TO_SIGNED(-463,11),
TO_SIGNED(-499,11),
TO_SIGNED(-533,11),
TO_SIGNED(-565,11),
TO_SIGNED(-595,11),
TO_SIGNED(-622,11),
TO_SIGNED(-647,11),
TO_SIGNED(-670,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-721,11),
TO_SIGNED(-733,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-720,11),
TO_SIGNED(-705,11),
TO_SIGNED(-688,11),
TO_SIGNED(-667,11),
TO_SIGNED(-645,11),
TO_SIGNED(-619,11),
TO_SIGNED(-592,11),
TO_SIGNED(-562,11),
TO_SIGNED(-529,11),
TO_SIGNED(-495,11),
TO_SIGNED(-459,11),
TO_SIGNED(-421,11),
TO_SIGNED(-381,11),
TO_SIGNED(-340,11),
TO_SIGNED(-297,11),
TO_SIGNED(-254,11),
TO_SIGNED(-209,11),
TO_SIGNED(-163,11),
TO_SIGNED(-117,11),
TO_SIGNED(-70,11),
TO_SIGNED(-24,11),
TO_SIGNED(24,11),
TO_SIGNED(70,11),
TO_SIGNED(117,11),
TO_SIGNED(163,11),
TO_SIGNED(209,11),
TO_SIGNED(254,11),
TO_SIGNED(297,11),
TO_SIGNED(340,11),
TO_SIGNED(381,11),
TO_SIGNED(421,11),
TO_SIGNED(459,11),
TO_SIGNED(495,11),
TO_SIGNED(529,11),
TO_SIGNED(562,11),
TO_SIGNED(592,11),
TO_SIGNED(619,11),
TO_SIGNED(645,11),
TO_SIGNED(667,11),
TO_SIGNED(688,11),
TO_SIGNED(705,11),
TO_SIGNED(720,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(733,11),
TO_SIGNED(721,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(670,11),
TO_SIGNED(647,11),
TO_SIGNED(622,11),
TO_SIGNED(595,11),
TO_SIGNED(565,11),
TO_SIGNED(533,11),
TO_SIGNED(499,11),
TO_SIGNED(463,11),
TO_SIGNED(425,11),
TO_SIGNED(386,11),
TO_SIGNED(345,11),
TO_SIGNED(302,11),
TO_SIGNED(259,11),
TO_SIGNED(214,11),
TO_SIGNED(168,11),
TO_SIGNED(122,11),
TO_SIGNED(76,11),
TO_SIGNED(29,11),
TO_SIGNED(-18,11),
TO_SIGNED(-65,11),
TO_SIGNED(-112,11),
TO_SIGNED(-158,11),
TO_SIGNED(-204,11),
TO_SIGNED(-248,11),
TO_SIGNED(-292,11),
TO_SIGNED(-335,11),
TO_SIGNED(-376,11),
TO_SIGNED(-416,11),
TO_SIGNED(-455,11),
TO_SIGNED(-491,11),
TO_SIGNED(-526,11),
TO_SIGNED(-558,11),
TO_SIGNED(-588,11),
TO_SIGNED(-616,11),
TO_SIGNED(-642,11),
TO_SIGNED(-665,11),
TO_SIGNED(-685,11),
TO_SIGNED(-703,11),
TO_SIGNED(-718,11),
TO_SIGNED(-730,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-692,11),
TO_SIGNED(-672,11),
TO_SIGNED(-650,11),
TO_SIGNED(-625,11),
TO_SIGNED(-598,11),
TO_SIGNED(-569,11),
TO_SIGNED(-537,11),
TO_SIGNED(-503,11),
TO_SIGNED(-467,11),
TO_SIGNED(-430,11),
TO_SIGNED(-390,11),
TO_SIGNED(-349,11),
TO_SIGNED(-307,11),
TO_SIGNED(-264,11),
TO_SIGNED(-219,11),
TO_SIGNED(-174,11),
TO_SIGNED(-128,11),
TO_SIGNED(-81,11),
TO_SIGNED(-34,11),
TO_SIGNED(13,11),
TO_SIGNED(60,11),
TO_SIGNED(106,11),
TO_SIGNED(153,11),
TO_SIGNED(198,11),
TO_SIGNED(243,11),
TO_SIGNED(287,11),
TO_SIGNED(330,11),
TO_SIGNED(372,11),
TO_SIGNED(412,11),
TO_SIGNED(450,11),
TO_SIGNED(487,11),
TO_SIGNED(522,11),
TO_SIGNED(554,11),
TO_SIGNED(585,11),
TO_SIGNED(613,11),
TO_SIGNED(639,11),
TO_SIGNED(662,11),
TO_SIGNED(683,11),
TO_SIGNED(701,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(724,11),
TO_SIGNED(710,11),
TO_SIGNED(694,11),
TO_SIGNED(675,11),
TO_SIGNED(653,11),
TO_SIGNED(628,11),
TO_SIGNED(601,11),
TO_SIGNED(572,11),
TO_SIGNED(541,11),
TO_SIGNED(507,11),
TO_SIGNED(471,11),
TO_SIGNED(434,11),
TO_SIGNED(395,11),
TO_SIGNED(354,11),
TO_SIGNED(312,11),
TO_SIGNED(269,11),
TO_SIGNED(224,11),
TO_SIGNED(179,11),
TO_SIGNED(133,11),
TO_SIGNED(86,11),
TO_SIGNED(40,11),
TO_SIGNED(-7,11),
TO_SIGNED(-54,11),
TO_SIGNED(-101,11),
TO_SIGNED(-148,11),
TO_SIGNED(-193,11),
TO_SIGNED(-238,11),
TO_SIGNED(-282,11),
TO_SIGNED(-325,11),
TO_SIGNED(-367,11),
TO_SIGNED(-407,11),
TO_SIGNED(-446,11),
TO_SIGNED(-483,11),
TO_SIGNED(-518,11),
TO_SIGNED(-551,11),
TO_SIGNED(-582,11),
TO_SIGNED(-610,11),
TO_SIGNED(-636,11),
TO_SIGNED(-660,11),
TO_SIGNED(-681,11),
TO_SIGNED(-699,11),
TO_SIGNED(-715,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-736,11),
TO_SIGNED(-725,11),
TO_SIGNED(-712,11),
TO_SIGNED(-696,11),
TO_SIGNED(-677,11),
TO_SIGNED(-655,11),
TO_SIGNED(-631,11),
TO_SIGNED(-605,11),
TO_SIGNED(-576,11),
TO_SIGNED(-544,11),
TO_SIGNED(-511,11),
TO_SIGNED(-476,11),
TO_SIGNED(-438,11),
TO_SIGNED(-399,11),
TO_SIGNED(-359,11),
TO_SIGNED(-317,11),
TO_SIGNED(-274,11),
TO_SIGNED(-229,11),
TO_SIGNED(-184,11),
TO_SIGNED(-138,11),
TO_SIGNED(-92,11),
TO_SIGNED(-45,11),
TO_SIGNED(2,11),
TO_SIGNED(49,11),
TO_SIGNED(96,11),
TO_SIGNED(142,11),
TO_SIGNED(188,11),
TO_SIGNED(233,11),
TO_SIGNED(277,11),
TO_SIGNED(321,11),
TO_SIGNED(362,11),
TO_SIGNED(403,11),
TO_SIGNED(442,11),
TO_SIGNED(479,11),
TO_SIGNED(514,11),
TO_SIGNED(547,11),
TO_SIGNED(578,11),
TO_SIGNED(607,11),
TO_SIGNED(633,11),
TO_SIGNED(657,11),
TO_SIGNED(679,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(698,11),
TO_SIGNED(679,11),
TO_SIGNED(658,11),
TO_SIGNED(634,11),
TO_SIGNED(608,11),
TO_SIGNED(579,11),
TO_SIGNED(548,11),
TO_SIGNED(515,11),
TO_SIGNED(480,11),
TO_SIGNED(443,11),
TO_SIGNED(404,11),
TO_SIGNED(363,11),
TO_SIGNED(322,11),
TO_SIGNED(278,11),
TO_SIGNED(234,11),
TO_SIGNED(189,11),
TO_SIGNED(143,11),
TO_SIGNED(97,11),
TO_SIGNED(50,11),
TO_SIGNED(3,11),
TO_SIGNED(-44,11),
TO_SIGNED(-91,11),
TO_SIGNED(-137,11),
TO_SIGNED(-183,11),
TO_SIGNED(-228,11),
TO_SIGNED(-273,11),
TO_SIGNED(-316,11),
TO_SIGNED(-358,11),
TO_SIGNED(-398,11),
TO_SIGNED(-437,11),
TO_SIGNED(-475,11),
TO_SIGNED(-510,11),
TO_SIGNED(-544,11),
TO_SIGNED(-575,11),
TO_SIGNED(-604,11),
TO_SIGNED(-631,11),
TO_SIGNED(-655,11),
TO_SIGNED(-676,11),
TO_SIGNED(-695,11),
TO_SIGNED(-712,11),
TO_SIGNED(-725,11),
TO_SIGNED(-736,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-715,11),
TO_SIGNED(-700,11),
TO_SIGNED(-681,11),
TO_SIGNED(-660,11),
TO_SIGNED(-637,11),
TO_SIGNED(-611,11),
TO_SIGNED(-582,11),
TO_SIGNED(-552,11),
TO_SIGNED(-519,11),
TO_SIGNED(-484,11),
TO_SIGNED(-447,11),
TO_SIGNED(-408,11),
TO_SIGNED(-368,11),
TO_SIGNED(-326,11),
TO_SIGNED(-283,11),
TO_SIGNED(-239,11),
TO_SIGNED(-194,11),
TO_SIGNED(-149,11),
TO_SIGNED(-102,11),
TO_SIGNED(-56,11),
TO_SIGNED(-9,11),
TO_SIGNED(38,11),
TO_SIGNED(85,11),
TO_SIGNED(132,11),
TO_SIGNED(178,11),
TO_SIGNED(223,11),
TO_SIGNED(268,11),
TO_SIGNED(311,11),
TO_SIGNED(353,11),
TO_SIGNED(394,11),
TO_SIGNED(433,11),
TO_SIGNED(471,11),
TO_SIGNED(506,11),
TO_SIGNED(540,11),
TO_SIGNED(571,11),
TO_SIGNED(601,11),
TO_SIGNED(628,11),
TO_SIGNED(652,11),
TO_SIGNED(674,11),
TO_SIGNED(693,11),
TO_SIGNED(710,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(739,11),
TO_SIGNED(729,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(684,11),
TO_SIGNED(663,11),
TO_SIGNED(640,11),
TO_SIGNED(614,11),
TO_SIGNED(586,11),
TO_SIGNED(555,11),
TO_SIGNED(523,11),
TO_SIGNED(488,11),
TO_SIGNED(451,11),
TO_SIGNED(413,11),
TO_SIGNED(373,11),
TO_SIGNED(331,11),
TO_SIGNED(288,11),
TO_SIGNED(244,11),
TO_SIGNED(200,11),
TO_SIGNED(154,11),
TO_SIGNED(108,11),
TO_SIGNED(61,11),
TO_SIGNED(14,11),
TO_SIGNED(-33,11),
TO_SIGNED(-80,11),
TO_SIGNED(-127,11),
TO_SIGNED(-173,11),
TO_SIGNED(-218,11),
TO_SIGNED(-263,11),
TO_SIGNED(-306,11),
TO_SIGNED(-348,11),
TO_SIGNED(-389,11),
TO_SIGNED(-429,11),
TO_SIGNED(-466,11),
TO_SIGNED(-502,11),
TO_SIGNED(-536,11),
TO_SIGNED(-568,11),
TO_SIGNED(-598,11),
TO_SIGNED(-625,11),
TO_SIGNED(-650,11),
TO_SIGNED(-672,11),
TO_SIGNED(-691,11),
TO_SIGNED(-708,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-686,11),
TO_SIGNED(-665,11),
TO_SIGNED(-642,11),
TO_SIGNED(-617,11),
TO_SIGNED(-589,11),
TO_SIGNED(-559,11),
TO_SIGNED(-526,11),
TO_SIGNED(-492,11),
TO_SIGNED(-455,11),
TO_SIGNED(-417,11),
TO_SIGNED(-377,11),
TO_SIGNED(-336,11),
TO_SIGNED(-293,11),
TO_SIGNED(-249,11),
TO_SIGNED(-205,11),
TO_SIGNED(-159,11),
TO_SIGNED(-113,11),
TO_SIGNED(-66,11),
TO_SIGNED(-19,11),
TO_SIGNED(28,11),
TO_SIGNED(75,11),
TO_SIGNED(121,11),
TO_SIGNED(167,11),
TO_SIGNED(213,11),
TO_SIGNED(258,11),
TO_SIGNED(301,11),
TO_SIGNED(344,11),
TO_SIGNED(385,11),
TO_SIGNED(424,11),
TO_SIGNED(462,11),
TO_SIGNED(498,11),
TO_SIGNED(532,11),
TO_SIGNED(564,11),
TO_SIGNED(594,11),
TO_SIGNED(622,11),
TO_SIGNED(647,11),
TO_SIGNED(669,11),
TO_SIGNED(689,11),
TO_SIGNED(706,11),
TO_SIGNED(721,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(720,11),
TO_SIGNED(705,11),
TO_SIGNED(688,11),
TO_SIGNED(668,11),
TO_SIGNED(645,11),
TO_SIGNED(620,11),
TO_SIGNED(592,11),
TO_SIGNED(562,11),
TO_SIGNED(530,11),
TO_SIGNED(496,11),
TO_SIGNED(460,11),
TO_SIGNED(422,11),
TO_SIGNED(382,11),
TO_SIGNED(341,11),
TO_SIGNED(298,11),
TO_SIGNED(255,11),
TO_SIGNED(210,11),
TO_SIGNED(164,11),
TO_SIGNED(118,11),
TO_SIGNED(71,11),
TO_SIGNED(25,11),
TO_SIGNED(-22,11),
TO_SIGNED(-69,11),
TO_SIGNED(-116,11),
TO_SIGNED(-162,11),
TO_SIGNED(-208,11),
TO_SIGNED(-252,11),
TO_SIGNED(-296,11),
TO_SIGNED(-339,11),
TO_SIGNED(-380,11),
TO_SIGNED(-420,11),
TO_SIGNED(-458,11),
TO_SIGNED(-494,11),
TO_SIGNED(-529,11),
TO_SIGNED(-561,11),
TO_SIGNED(-591,11),
TO_SIGNED(-619,11),
TO_SIGNED(-644,11),
TO_SIGNED(-667,11),
TO_SIGNED(-687,11),
TO_SIGNED(-705,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-733,11),
TO_SIGNED(-721,11),
TO_SIGNED(-707,11),
TO_SIGNED(-690,11),
TO_SIGNED(-670,11),
TO_SIGNED(-648,11),
TO_SIGNED(-623,11),
TO_SIGNED(-596,11),
TO_SIGNED(-566,11),
TO_SIGNED(-534,11),
TO_SIGNED(-500,11),
TO_SIGNED(-464,11),
TO_SIGNED(-426,11),
TO_SIGNED(-387,11),
TO_SIGNED(-345,11),
TO_SIGNED(-303,11),
TO_SIGNED(-260,11),
TO_SIGNED(-215,11),
TO_SIGNED(-169,11),
TO_SIGNED(-123,11),
TO_SIGNED(-77,11),
TO_SIGNED(-30,11),
TO_SIGNED(17,11),
TO_SIGNED(64,11),
TO_SIGNED(111,11),
TO_SIGNED(157,11),
TO_SIGNED(203,11),
TO_SIGNED(247,11),
TO_SIGNED(291,11),
TO_SIGNED(334,11),
TO_SIGNED(375,11),
TO_SIGNED(415,11),
TO_SIGNED(454,11),
TO_SIGNED(490,11),
TO_SIGNED(525,11),
TO_SIGNED(557,11),
TO_SIGNED(588,11),
TO_SIGNED(616,11),
TO_SIGNED(641,11),
TO_SIGNED(664,11),
TO_SIGNED(685,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(709,11),
TO_SIGNED(692,11),
TO_SIGNED(673,11),
TO_SIGNED(651,11),
TO_SIGNED(626,11),
TO_SIGNED(599,11),
TO_SIGNED(569,11),
TO_SIGNED(538,11),
TO_SIGNED(504,11),
TO_SIGNED(468,11),
TO_SIGNED(430,11),
TO_SIGNED(391,11),
TO_SIGNED(350,11),
TO_SIGNED(308,11),
TO_SIGNED(265,11),
TO_SIGNED(220,11),
TO_SIGNED(175,11),
TO_SIGNED(129,11),
TO_SIGNED(82,11),
TO_SIGNED(35,11),
TO_SIGNED(-12,11),
TO_SIGNED(-59,11),
TO_SIGNED(-105,11),
TO_SIGNED(-152,11),
TO_SIGNED(-197,11),
TO_SIGNED(-242,11),
TO_SIGNED(-286,11),
TO_SIGNED(-329,11),
TO_SIGNED(-371,11),
TO_SIGNED(-411,11),
TO_SIGNED(-449,11),
TO_SIGNED(-486,11),
TO_SIGNED(-521,11),
TO_SIGNED(-554,11),
TO_SIGNED(-584,11),
TO_SIGNED(-613,11),
TO_SIGNED(-639,11),
TO_SIGNED(-662,11),
TO_SIGNED(-683,11),
TO_SIGNED(-701,11),
TO_SIGNED(-716,11),
TO_SIGNED(-729,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-711,11),
TO_SIGNED(-694,11),
TO_SIGNED(-675,11),
TO_SIGNED(-653,11),
TO_SIGNED(-629,11),
TO_SIGNED(-602,11),
TO_SIGNED(-573,11),
TO_SIGNED(-541,11),
TO_SIGNED(-508,11),
TO_SIGNED(-472,11),
TO_SIGNED(-435,11),
TO_SIGNED(-396,11),
TO_SIGNED(-355,11),
TO_SIGNED(-313,11),
TO_SIGNED(-270,11),
TO_SIGNED(-225,11),
TO_SIGNED(-180,11),
TO_SIGNED(-134,11),
TO_SIGNED(-87,11),
TO_SIGNED(-41,11),
TO_SIGNED(6,11),
TO_SIGNED(53,11),
TO_SIGNED(100,11),
TO_SIGNED(147,11),
TO_SIGNED(192,11),
TO_SIGNED(237,11),
TO_SIGNED(281,11),
TO_SIGNED(324,11),
TO_SIGNED(366,11),
TO_SIGNED(406,11),
TO_SIGNED(445,11),
TO_SIGNED(482,11),
TO_SIGNED(517,11),
TO_SIGNED(550,11),
TO_SIGNED(581,11),
TO_SIGNED(610,11),
TO_SIGNED(636,11),
TO_SIGNED(659,11),
TO_SIGNED(681,11),
TO_SIGNED(699,11),
TO_SIGNED(715,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(712,11),
TO_SIGNED(696,11),
TO_SIGNED(677,11),
TO_SIGNED(656,11),
TO_SIGNED(632,11),
TO_SIGNED(605,11),
TO_SIGNED(576,11),
TO_SIGNED(545,11),
TO_SIGNED(512,11),
TO_SIGNED(476,11),
TO_SIGNED(439,11),
TO_SIGNED(400,11),
TO_SIGNED(360,11),
TO_SIGNED(318,11),
TO_SIGNED(275,11),
TO_SIGNED(230,11),
TO_SIGNED(185,11),
TO_SIGNED(139,11),
TO_SIGNED(93,11),
TO_SIGNED(46,11),
TO_SIGNED(-1,11),
TO_SIGNED(-48,11),
TO_SIGNED(-95,11),
TO_SIGNED(-141,11),
TO_SIGNED(-187,11),
TO_SIGNED(-232,11),
TO_SIGNED(-276,11),
TO_SIGNED(-320,11),
TO_SIGNED(-362,11),
TO_SIGNED(-402,11),
TO_SIGNED(-441,11),
TO_SIGNED(-478,11),
TO_SIGNED(-513,11),
TO_SIGNED(-547,11),
TO_SIGNED(-578,11),
TO_SIGNED(-606,11),
TO_SIGNED(-633,11),
TO_SIGNED(-657,11),
TO_SIGNED(-678,11),
TO_SIGNED(-697,11),
TO_SIGNED(-713,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-714,11),
TO_SIGNED(-698,11),
TO_SIGNED(-680,11),
TO_SIGNED(-658,11),
TO_SIGNED(-635,11),
TO_SIGNED(-608,11),
TO_SIGNED(-580,11),
TO_SIGNED(-549,11),
TO_SIGNED(-516,11),
TO_SIGNED(-480,11),
TO_SIGNED(-443,11),
TO_SIGNED(-405,11),
TO_SIGNED(-364,11),
TO_SIGNED(-323,11),
TO_SIGNED(-279,11),
TO_SIGNED(-235,11),
TO_SIGNED(-190,11),
TO_SIGNED(-144,11),
TO_SIGNED(-98,11),
TO_SIGNED(-51,11),
TO_SIGNED(-4,11),
TO_SIGNED(43,11),
TO_SIGNED(90,11),
TO_SIGNED(136,11),
TO_SIGNED(182,11),
TO_SIGNED(227,11),
TO_SIGNED(272,11),
TO_SIGNED(315,11),
TO_SIGNED(357,11),
TO_SIGNED(397,11),
TO_SIGNED(437,11),
TO_SIGNED(474,11),
TO_SIGNED(509,11),
TO_SIGNED(543,11),
TO_SIGNED(574,11),
TO_SIGNED(603,11),
TO_SIGNED(630,11),
TO_SIGNED(654,11),
TO_SIGNED(676,11),
TO_SIGNED(695,11),
TO_SIGNED(711,11),
TO_SIGNED(725,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(716,11),
TO_SIGNED(700,11),
TO_SIGNED(682,11),
TO_SIGNED(661,11),
TO_SIGNED(637,11),
TO_SIGNED(611,11),
TO_SIGNED(583,11),
TO_SIGNED(552,11),
TO_SIGNED(519,11),
TO_SIGNED(485,11),
TO_SIGNED(448,11),
TO_SIGNED(409,11),
TO_SIGNED(369,11),
TO_SIGNED(327,11),
TO_SIGNED(284,11),
TO_SIGNED(240,11),
TO_SIGNED(195,11),
TO_SIGNED(150,11),
TO_SIGNED(103,11),
TO_SIGNED(57,11),
TO_SIGNED(10,11),
TO_SIGNED(-37,11),
TO_SIGNED(-84,11),
TO_SIGNED(-131,11),
TO_SIGNED(-177,11),
TO_SIGNED(-222,11),
TO_SIGNED(-267,11),
TO_SIGNED(-310,11),
TO_SIGNED(-352,11),
TO_SIGNED(-393,11),
TO_SIGNED(-432,11),
TO_SIGNED(-470,11),
TO_SIGNED(-505,11),
TO_SIGNED(-539,11),
TO_SIGNED(-571,11),
TO_SIGNED(-600,11),
TO_SIGNED(-627,11),
TO_SIGNED(-652,11),
TO_SIGNED(-674,11),
TO_SIGNED(-693,11),
TO_SIGNED(-710,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-702,11),
TO_SIGNED(-684,11),
TO_SIGNED(-663,11),
TO_SIGNED(-640,11),
TO_SIGNED(-615,11),
TO_SIGNED(-586,11),
TO_SIGNED(-556,11),
TO_SIGNED(-523,11),
TO_SIGNED(-489,11),
TO_SIGNED(-452,11),
TO_SIGNED(-414,11),
TO_SIGNED(-374,11),
TO_SIGNED(-332,11),
TO_SIGNED(-289,11),
TO_SIGNED(-245,11),
TO_SIGNED(-201,11),
TO_SIGNED(-155,11),
TO_SIGNED(-109,11),
TO_SIGNED(-62,11),
TO_SIGNED(-15,11),
TO_SIGNED(32,11),
TO_SIGNED(79,11),
TO_SIGNED(125,11),
TO_SIGNED(172,11),
TO_SIGNED(217,11),
TO_SIGNED(262,11),
TO_SIGNED(305,11),
TO_SIGNED(347,11),
TO_SIGNED(388,11),
TO_SIGNED(428,11),
TO_SIGNED(466,11),
TO_SIGNED(501,11),
TO_SIGNED(535,11),
TO_SIGNED(567,11),
TO_SIGNED(597,11),
TO_SIGNED(624,11),
TO_SIGNED(649,11),
TO_SIGNED(671,11),
TO_SIGNED(691,11),
TO_SIGNED(708,11),
TO_SIGNED(722,11),
TO_SIGNED(733,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(704,11),
TO_SIGNED(686,11),
TO_SIGNED(666,11),
TO_SIGNED(643,11),
TO_SIGNED(618,11),
TO_SIGNED(590,11),
TO_SIGNED(559,11),
TO_SIGNED(527,11),
TO_SIGNED(493,11),
TO_SIGNED(456,11),
TO_SIGNED(418,11),
TO_SIGNED(378,11),
TO_SIGNED(337,11),
TO_SIGNED(294,11),
TO_SIGNED(250,11),
TO_SIGNED(206,11),
TO_SIGNED(160,11),
TO_SIGNED(114,11),
TO_SIGNED(67,11),
TO_SIGNED(20,11),
TO_SIGNED(-27,11),
TO_SIGNED(-74,11),
TO_SIGNED(-120,11),
TO_SIGNED(-166,11),
TO_SIGNED(-212,11),
TO_SIGNED(-257,11),
TO_SIGNED(-300,11),
TO_SIGNED(-343,11),
TO_SIGNED(-384,11),
TO_SIGNED(-423,11),
TO_SIGNED(-461,11),
TO_SIGNED(-497,11),
TO_SIGNED(-532,11),
TO_SIGNED(-564,11),
TO_SIGNED(-594,11),
TO_SIGNED(-621,11),
TO_SIGNED(-646,11),
TO_SIGNED(-669,11),
TO_SIGNED(-689,11),
TO_SIGNED(-706,11),
TO_SIGNED(-721,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-720,11),
TO_SIGNED(-706,11),
TO_SIGNED(-688,11),
TO_SIGNED(-668,11),
TO_SIGNED(-646,11),
TO_SIGNED(-621,11),
TO_SIGNED(-593,11),
TO_SIGNED(-563,11),
TO_SIGNED(-531,11),
TO_SIGNED(-497,11),
TO_SIGNED(-460,11),
TO_SIGNED(-422,11),
TO_SIGNED(-383,11),
TO_SIGNED(-342,11),
TO_SIGNED(-299,11),
TO_SIGNED(-256,11),
TO_SIGNED(-211,11),
TO_SIGNED(-165,11),
TO_SIGNED(-119,11),
TO_SIGNED(-73,11),
TO_SIGNED(-26,11),
TO_SIGNED(21,11),
TO_SIGNED(68,11),
TO_SIGNED(115,11),
TO_SIGNED(161,11),
TO_SIGNED(207,11),
TO_SIGNED(251,11),
TO_SIGNED(295,11),
TO_SIGNED(338,11),
TO_SIGNED(379,11),
TO_SIGNED(419,11),
TO_SIGNED(457,11),
TO_SIGNED(493,11),
TO_SIGNED(528,11),
TO_SIGNED(560,11),
TO_SIGNED(590,11),
TO_SIGNED(618,11),
TO_SIGNED(644,11),
TO_SIGNED(666,11),
TO_SIGNED(687,11),
TO_SIGNED(704,11),
TO_SIGNED(719,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(671,11),
TO_SIGNED(648,11),
TO_SIGNED(624,11),
TO_SIGNED(596,11),
TO_SIGNED(567,11),
TO_SIGNED(535,11),
TO_SIGNED(501,11),
TO_SIGNED(465,11),
TO_SIGNED(427,11),
TO_SIGNED(387,11),
TO_SIGNED(346,11),
TO_SIGNED(304,11),
TO_SIGNED(261,11),
TO_SIGNED(216,11),
TO_SIGNED(171,11),
TO_SIGNED(124,11),
TO_SIGNED(78,11),
TO_SIGNED(31,11),
TO_SIGNED(-16,11),
TO_SIGNED(-63,11),
TO_SIGNED(-110,11),
TO_SIGNED(-156,11),
TO_SIGNED(-202,11),
TO_SIGNED(-246,11),
TO_SIGNED(-290,11),
TO_SIGNED(-333,11),
TO_SIGNED(-375,11),
TO_SIGNED(-415,11),
TO_SIGNED(-453,11),
TO_SIGNED(-489,11),
TO_SIGNED(-524,11),
TO_SIGNED(-557,11),
TO_SIGNED(-587,11),
TO_SIGNED(-615,11),
TO_SIGNED(-641,11),
TO_SIGNED(-664,11),
TO_SIGNED(-685,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-730,11),
TO_SIGNED(-739,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-693,11),
TO_SIGNED(-673,11),
TO_SIGNED(-651,11),
TO_SIGNED(-627,11),
TO_SIGNED(-599,11),
TO_SIGNED(-570,11),
TO_SIGNED(-538,11),
TO_SIGNED(-505,11),
TO_SIGNED(-469,11),
TO_SIGNED(-431,11),
TO_SIGNED(-392,11),
TO_SIGNED(-351,11),
TO_SIGNED(-309,11),
TO_SIGNED(-266,11),
TO_SIGNED(-221,11),
TO_SIGNED(-176,11),
TO_SIGNED(-130,11),
TO_SIGNED(-83,11),
TO_SIGNED(-36,11),
TO_SIGNED(11,11),
TO_SIGNED(58,11),
TO_SIGNED(104,11),
TO_SIGNED(151,11),
TO_SIGNED(196,11),
TO_SIGNED(241,11),
TO_SIGNED(285,11),
TO_SIGNED(328,11),
TO_SIGNED(370,11),
TO_SIGNED(410,11),
TO_SIGNED(449,11),
TO_SIGNED(485,11),
TO_SIGNED(520,11),
TO_SIGNED(553,11),
TO_SIGNED(584,11),
TO_SIGNED(612,11),
TO_SIGNED(638,11),
TO_SIGNED(661,11),
TO_SIGNED(682,11),
TO_SIGNED(700,11),
TO_SIGNED(716,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(725,11),
TO_SIGNED(711,11),
TO_SIGNED(695,11),
TO_SIGNED(675,11),
TO_SIGNED(654,11),
TO_SIGNED(629,11),
TO_SIGNED(603,11),
TO_SIGNED(574,11),
TO_SIGNED(542,11),
TO_SIGNED(509,11),
TO_SIGNED(473,11),
TO_SIGNED(436,11),
TO_SIGNED(397,11),
TO_SIGNED(356,11),
TO_SIGNED(314,11),
TO_SIGNED(271,11),
TO_SIGNED(226,11),
TO_SIGNED(181,11),
TO_SIGNED(135,11),
TO_SIGNED(88,11),
TO_SIGNED(42,11),
TO_SIGNED(-5,11),
TO_SIGNED(-52,11),
TO_SIGNED(-99,11),
TO_SIGNED(-145,11),
TO_SIGNED(-191,11),
TO_SIGNED(-236,11),
TO_SIGNED(-280,11),
TO_SIGNED(-323,11),
TO_SIGNED(-365,11),
TO_SIGNED(-406,11),
TO_SIGNED(-444,11),
TO_SIGNED(-481,11),
TO_SIGNED(-516,11),
TO_SIGNED(-549,11),
TO_SIGNED(-580,11),
TO_SIGNED(-609,11),
TO_SIGNED(-635,11),
TO_SIGNED(-659,11),
TO_SIGNED(-680,11),
TO_SIGNED(-699,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-736,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-678,11),
TO_SIGNED(-656,11),
TO_SIGNED(-632,11),
TO_SIGNED(-606,11),
TO_SIGNED(-577,11),
TO_SIGNED(-546,11),
TO_SIGNED(-512,11),
TO_SIGNED(-477,11),
TO_SIGNED(-440,11),
TO_SIGNED(-401,11),
TO_SIGNED(-361,11),
TO_SIGNED(-319,11),
TO_SIGNED(-275,11),
TO_SIGNED(-231,11),
TO_SIGNED(-186,11),
TO_SIGNED(-140,11),
TO_SIGNED(-94,11),
TO_SIGNED(-47,11),
TO_SIGNED(0,11),
TO_SIGNED(47,11),
TO_SIGNED(94,11),
TO_SIGNED(140,11),
TO_SIGNED(186,11),
TO_SIGNED(231,11),
TO_SIGNED(275,11),
TO_SIGNED(319,11),
TO_SIGNED(361,11),
TO_SIGNED(401,11),
TO_SIGNED(440,11),
TO_SIGNED(477,11),
TO_SIGNED(512,11),
TO_SIGNED(546,11),
TO_SIGNED(577,11),
TO_SIGNED(606,11),
TO_SIGNED(632,11),
TO_SIGNED(656,11),
TO_SIGNED(678,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(736,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(699,11),
TO_SIGNED(680,11),
TO_SIGNED(659,11),
TO_SIGNED(635,11),
TO_SIGNED(609,11),
TO_SIGNED(580,11),
TO_SIGNED(549,11),
TO_SIGNED(516,11),
TO_SIGNED(481,11),
TO_SIGNED(444,11),
TO_SIGNED(406,11),
TO_SIGNED(365,11),
TO_SIGNED(323,11),
TO_SIGNED(280,11),
TO_SIGNED(236,11),
TO_SIGNED(191,11),
TO_SIGNED(145,11),
TO_SIGNED(99,11),
TO_SIGNED(52,11),
TO_SIGNED(5,11),
TO_SIGNED(-42,11),
TO_SIGNED(-88,11),
TO_SIGNED(-135,11),
TO_SIGNED(-181,11),
TO_SIGNED(-226,11),
TO_SIGNED(-271,11),
TO_SIGNED(-314,11),
TO_SIGNED(-356,11),
TO_SIGNED(-397,11),
TO_SIGNED(-436,11),
TO_SIGNED(-473,11),
TO_SIGNED(-509,11),
TO_SIGNED(-542,11),
TO_SIGNED(-574,11),
TO_SIGNED(-603,11),
TO_SIGNED(-629,11),
TO_SIGNED(-654,11),
TO_SIGNED(-675,11),
TO_SIGNED(-695,11),
TO_SIGNED(-711,11),
TO_SIGNED(-725,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-716,11),
TO_SIGNED(-700,11),
TO_SIGNED(-682,11),
TO_SIGNED(-661,11),
TO_SIGNED(-638,11),
TO_SIGNED(-612,11),
TO_SIGNED(-584,11),
TO_SIGNED(-553,11),
TO_SIGNED(-520,11),
TO_SIGNED(-485,11),
TO_SIGNED(-449,11),
TO_SIGNED(-410,11),
TO_SIGNED(-370,11),
TO_SIGNED(-328,11),
TO_SIGNED(-285,11),
TO_SIGNED(-241,11),
TO_SIGNED(-196,11),
TO_SIGNED(-151,11),
TO_SIGNED(-104,11),
TO_SIGNED(-58,11),
TO_SIGNED(-11,11),
TO_SIGNED(36,11),
TO_SIGNED(83,11),
TO_SIGNED(130,11),
TO_SIGNED(176,11),
TO_SIGNED(221,11),
TO_SIGNED(266,11),
TO_SIGNED(309,11),
TO_SIGNED(351,11),
TO_SIGNED(392,11),
TO_SIGNED(431,11),
TO_SIGNED(469,11),
TO_SIGNED(505,11),
TO_SIGNED(538,11),
TO_SIGNED(570,11),
TO_SIGNED(599,11),
TO_SIGNED(627,11),
TO_SIGNED(651,11),
TO_SIGNED(673,11),
TO_SIGNED(693,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(739,11),
TO_SIGNED(730,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(685,11),
TO_SIGNED(664,11),
TO_SIGNED(641,11),
TO_SIGNED(615,11),
TO_SIGNED(587,11),
TO_SIGNED(557,11),
TO_SIGNED(524,11),
TO_SIGNED(489,11),
TO_SIGNED(453,11),
TO_SIGNED(415,11),
TO_SIGNED(375,11),
TO_SIGNED(333,11),
TO_SIGNED(290,11),
TO_SIGNED(246,11),
TO_SIGNED(202,11),
TO_SIGNED(156,11),
TO_SIGNED(110,11),
TO_SIGNED(63,11),
TO_SIGNED(16,11),
TO_SIGNED(-31,11),
TO_SIGNED(-78,11),
TO_SIGNED(-124,11),
TO_SIGNED(-171,11),
TO_SIGNED(-216,11),
TO_SIGNED(-261,11),
TO_SIGNED(-304,11),
TO_SIGNED(-346,11),
TO_SIGNED(-387,11),
TO_SIGNED(-427,11),
TO_SIGNED(-465,11),
TO_SIGNED(-501,11),
TO_SIGNED(-535,11),
TO_SIGNED(-567,11),
TO_SIGNED(-596,11),
TO_SIGNED(-624,11),
TO_SIGNED(-648,11),
TO_SIGNED(-671,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-719,11),
TO_SIGNED(-704,11),
TO_SIGNED(-687,11),
TO_SIGNED(-666,11),
TO_SIGNED(-644,11),
TO_SIGNED(-618,11),
TO_SIGNED(-590,11),
TO_SIGNED(-560,11),
TO_SIGNED(-528,11),
TO_SIGNED(-493,11),
TO_SIGNED(-457,11),
TO_SIGNED(-419,11),
TO_SIGNED(-379,11),
TO_SIGNED(-338,11),
TO_SIGNED(-295,11),
TO_SIGNED(-251,11),
TO_SIGNED(-207,11),
TO_SIGNED(-161,11),
TO_SIGNED(-115,11),
TO_SIGNED(-68,11),
TO_SIGNED(-21,11),
TO_SIGNED(26,11),
TO_SIGNED(73,11),
TO_SIGNED(119,11),
TO_SIGNED(165,11),
TO_SIGNED(211,11),
TO_SIGNED(256,11),
TO_SIGNED(299,11),
TO_SIGNED(342,11),
TO_SIGNED(383,11),
TO_SIGNED(422,11),
TO_SIGNED(460,11),
TO_SIGNED(497,11),
TO_SIGNED(531,11),
TO_SIGNED(563,11),
TO_SIGNED(593,11),
TO_SIGNED(621,11),
TO_SIGNED(646,11),
TO_SIGNED(668,11),
TO_SIGNED(688,11),
TO_SIGNED(706,11),
TO_SIGNED(720,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(721,11),
TO_SIGNED(706,11),
TO_SIGNED(689,11),
TO_SIGNED(669,11),
TO_SIGNED(646,11),
TO_SIGNED(621,11),
TO_SIGNED(594,11),
TO_SIGNED(564,11),
TO_SIGNED(532,11),
TO_SIGNED(497,11),
TO_SIGNED(461,11),
TO_SIGNED(423,11),
TO_SIGNED(384,11),
TO_SIGNED(343,11),
TO_SIGNED(300,11),
TO_SIGNED(257,11),
TO_SIGNED(212,11),
TO_SIGNED(166,11),
TO_SIGNED(120,11),
TO_SIGNED(74,11),
TO_SIGNED(27,11),
TO_SIGNED(-20,11),
TO_SIGNED(-67,11),
TO_SIGNED(-114,11),
TO_SIGNED(-160,11),
TO_SIGNED(-206,11),
TO_SIGNED(-250,11),
TO_SIGNED(-294,11),
TO_SIGNED(-337,11),
TO_SIGNED(-378,11),
TO_SIGNED(-418,11),
TO_SIGNED(-456,11),
TO_SIGNED(-493,11),
TO_SIGNED(-527,11),
TO_SIGNED(-559,11),
TO_SIGNED(-590,11),
TO_SIGNED(-618,11),
TO_SIGNED(-643,11),
TO_SIGNED(-666,11),
TO_SIGNED(-686,11),
TO_SIGNED(-704,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-733,11),
TO_SIGNED(-722,11),
TO_SIGNED(-708,11),
TO_SIGNED(-691,11),
TO_SIGNED(-671,11),
TO_SIGNED(-649,11),
TO_SIGNED(-624,11),
TO_SIGNED(-597,11),
TO_SIGNED(-567,11),
TO_SIGNED(-535,11),
TO_SIGNED(-501,11),
TO_SIGNED(-466,11),
TO_SIGNED(-428,11),
TO_SIGNED(-388,11),
TO_SIGNED(-347,11),
TO_SIGNED(-305,11),
TO_SIGNED(-262,11),
TO_SIGNED(-217,11),
TO_SIGNED(-172,11),
TO_SIGNED(-125,11),
TO_SIGNED(-79,11),
TO_SIGNED(-32,11),
TO_SIGNED(15,11),
TO_SIGNED(62,11),
TO_SIGNED(109,11),
TO_SIGNED(155,11),
TO_SIGNED(201,11),
TO_SIGNED(245,11),
TO_SIGNED(289,11),
TO_SIGNED(332,11),
TO_SIGNED(374,11),
TO_SIGNED(414,11),
TO_SIGNED(452,11),
TO_SIGNED(489,11),
TO_SIGNED(523,11),
TO_SIGNED(556,11),
TO_SIGNED(586,11),
TO_SIGNED(615,11),
TO_SIGNED(640,11),
TO_SIGNED(663,11),
TO_SIGNED(684,11),
TO_SIGNED(702,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(710,11),
TO_SIGNED(693,11),
TO_SIGNED(674,11),
TO_SIGNED(652,11),
TO_SIGNED(627,11),
TO_SIGNED(600,11),
TO_SIGNED(571,11),
TO_SIGNED(539,11),
TO_SIGNED(505,11),
TO_SIGNED(470,11),
TO_SIGNED(432,11),
TO_SIGNED(393,11),
TO_SIGNED(352,11),
TO_SIGNED(310,11),
TO_SIGNED(267,11),
TO_SIGNED(222,11),
TO_SIGNED(177,11),
TO_SIGNED(131,11),
TO_SIGNED(84,11),
TO_SIGNED(37,11),
TO_SIGNED(-10,11),
TO_SIGNED(-57,11),
TO_SIGNED(-103,11),
TO_SIGNED(-150,11),
TO_SIGNED(-195,11),
TO_SIGNED(-240,11),
TO_SIGNED(-284,11),
TO_SIGNED(-327,11),
TO_SIGNED(-369,11),
TO_SIGNED(-409,11),
TO_SIGNED(-448,11),
TO_SIGNED(-485,11),
TO_SIGNED(-519,11),
TO_SIGNED(-552,11),
TO_SIGNED(-583,11),
TO_SIGNED(-611,11),
TO_SIGNED(-637,11),
TO_SIGNED(-661,11),
TO_SIGNED(-682,11),
TO_SIGNED(-700,11),
TO_SIGNED(-716,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-725,11),
TO_SIGNED(-711,11),
TO_SIGNED(-695,11),
TO_SIGNED(-676,11),
TO_SIGNED(-654,11),
TO_SIGNED(-630,11),
TO_SIGNED(-603,11),
TO_SIGNED(-574,11),
TO_SIGNED(-543,11),
TO_SIGNED(-509,11),
TO_SIGNED(-474,11),
TO_SIGNED(-437,11),
TO_SIGNED(-397,11),
TO_SIGNED(-357,11),
TO_SIGNED(-315,11),
TO_SIGNED(-272,11),
TO_SIGNED(-227,11),
TO_SIGNED(-182,11),
TO_SIGNED(-136,11),
TO_SIGNED(-90,11),
TO_SIGNED(-43,11),
TO_SIGNED(4,11),
TO_SIGNED(51,11),
TO_SIGNED(98,11),
TO_SIGNED(144,11),
TO_SIGNED(190,11),
TO_SIGNED(235,11),
TO_SIGNED(279,11),
TO_SIGNED(323,11),
TO_SIGNED(364,11),
TO_SIGNED(405,11),
TO_SIGNED(443,11),
TO_SIGNED(480,11),
TO_SIGNED(516,11),
TO_SIGNED(549,11),
TO_SIGNED(580,11),
TO_SIGNED(608,11),
TO_SIGNED(635,11),
TO_SIGNED(658,11),
TO_SIGNED(680,11),
TO_SIGNED(698,11),
TO_SIGNED(714,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(713,11),
TO_SIGNED(697,11),
TO_SIGNED(678,11),
TO_SIGNED(657,11),
TO_SIGNED(633,11),
TO_SIGNED(606,11),
TO_SIGNED(578,11),
TO_SIGNED(547,11),
TO_SIGNED(513,11),
TO_SIGNED(478,11),
TO_SIGNED(441,11),
TO_SIGNED(402,11),
TO_SIGNED(362,11),
TO_SIGNED(320,11),
TO_SIGNED(276,11),
TO_SIGNED(232,11),
TO_SIGNED(187,11),
TO_SIGNED(141,11),
TO_SIGNED(95,11),
TO_SIGNED(48,11),
TO_SIGNED(1,11),
TO_SIGNED(-46,11),
TO_SIGNED(-93,11),
TO_SIGNED(-139,11),
TO_SIGNED(-185,11),
TO_SIGNED(-230,11),
TO_SIGNED(-275,11),
TO_SIGNED(-318,11),
TO_SIGNED(-360,11),
TO_SIGNED(-400,11),
TO_SIGNED(-439,11),
TO_SIGNED(-476,11),
TO_SIGNED(-512,11),
TO_SIGNED(-545,11),
TO_SIGNED(-576,11),
TO_SIGNED(-605,11),
TO_SIGNED(-632,11),
TO_SIGNED(-656,11),
TO_SIGNED(-677,11),
TO_SIGNED(-696,11),
TO_SIGNED(-712,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-715,11),
TO_SIGNED(-699,11),
TO_SIGNED(-681,11),
TO_SIGNED(-659,11),
TO_SIGNED(-636,11),
TO_SIGNED(-610,11),
TO_SIGNED(-581,11),
TO_SIGNED(-550,11),
TO_SIGNED(-517,11),
TO_SIGNED(-482,11),
TO_SIGNED(-445,11),
TO_SIGNED(-406,11),
TO_SIGNED(-366,11),
TO_SIGNED(-324,11),
TO_SIGNED(-281,11),
TO_SIGNED(-237,11),
TO_SIGNED(-192,11),
TO_SIGNED(-147,11),
TO_SIGNED(-100,11),
TO_SIGNED(-53,11),
TO_SIGNED(-6,11),
TO_SIGNED(41,11),
TO_SIGNED(87,11),
TO_SIGNED(134,11),
TO_SIGNED(180,11),
TO_SIGNED(225,11),
TO_SIGNED(270,11),
TO_SIGNED(313,11),
TO_SIGNED(355,11),
TO_SIGNED(396,11),
TO_SIGNED(435,11),
TO_SIGNED(472,11),
TO_SIGNED(508,11),
TO_SIGNED(541,11),
TO_SIGNED(573,11),
TO_SIGNED(602,11),
TO_SIGNED(629,11),
TO_SIGNED(653,11),
TO_SIGNED(675,11),
TO_SIGNED(694,11),
TO_SIGNED(711,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(729,11),
TO_SIGNED(716,11),
TO_SIGNED(701,11),
TO_SIGNED(683,11),
TO_SIGNED(662,11),
TO_SIGNED(639,11),
TO_SIGNED(613,11),
TO_SIGNED(584,11),
TO_SIGNED(554,11),
TO_SIGNED(521,11),
TO_SIGNED(486,11),
TO_SIGNED(449,11),
TO_SIGNED(411,11),
TO_SIGNED(371,11),
TO_SIGNED(329,11),
TO_SIGNED(286,11),
TO_SIGNED(242,11),
TO_SIGNED(197,11),
TO_SIGNED(152,11),
TO_SIGNED(105,11),
TO_SIGNED(59,11),
TO_SIGNED(12,11),
TO_SIGNED(-35,11),
TO_SIGNED(-82,11),
TO_SIGNED(-129,11),
TO_SIGNED(-175,11),
TO_SIGNED(-220,11),
TO_SIGNED(-265,11),
TO_SIGNED(-308,11),
TO_SIGNED(-350,11),
TO_SIGNED(-391,11),
TO_SIGNED(-430,11),
TO_SIGNED(-468,11),
TO_SIGNED(-504,11),
TO_SIGNED(-538,11),
TO_SIGNED(-569,11),
TO_SIGNED(-599,11),
TO_SIGNED(-626,11),
TO_SIGNED(-651,11),
TO_SIGNED(-673,11),
TO_SIGNED(-692,11),
TO_SIGNED(-709,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-685,11),
TO_SIGNED(-664,11),
TO_SIGNED(-641,11),
TO_SIGNED(-616,11),
TO_SIGNED(-588,11),
TO_SIGNED(-557,11),
TO_SIGNED(-525,11),
TO_SIGNED(-490,11),
TO_SIGNED(-454,11),
TO_SIGNED(-415,11),
TO_SIGNED(-375,11),
TO_SIGNED(-334,11),
TO_SIGNED(-291,11),
TO_SIGNED(-247,11),
TO_SIGNED(-203,11),
TO_SIGNED(-157,11),
TO_SIGNED(-111,11),
TO_SIGNED(-64,11),
TO_SIGNED(-17,11),
TO_SIGNED(30,11),
TO_SIGNED(77,11),
TO_SIGNED(123,11),
TO_SIGNED(169,11),
TO_SIGNED(215,11),
TO_SIGNED(260,11),
TO_SIGNED(303,11),
TO_SIGNED(345,11),
TO_SIGNED(387,11),
TO_SIGNED(426,11),
TO_SIGNED(464,11),
TO_SIGNED(500,11),
TO_SIGNED(534,11),
TO_SIGNED(566,11),
TO_SIGNED(596,11),
TO_SIGNED(623,11),
TO_SIGNED(648,11),
TO_SIGNED(670,11),
TO_SIGNED(690,11),
TO_SIGNED(707,11),
TO_SIGNED(721,11),
TO_SIGNED(733,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(705,11),
TO_SIGNED(687,11),
TO_SIGNED(667,11),
TO_SIGNED(644,11),
TO_SIGNED(619,11),
TO_SIGNED(591,11),
TO_SIGNED(561,11),
TO_SIGNED(529,11),
TO_SIGNED(494,11),
TO_SIGNED(458,11),
TO_SIGNED(420,11),
TO_SIGNED(380,11),
TO_SIGNED(339,11),
TO_SIGNED(296,11),
TO_SIGNED(252,11),
TO_SIGNED(208,11),
TO_SIGNED(162,11),
TO_SIGNED(116,11),
TO_SIGNED(69,11),
TO_SIGNED(22,11),
TO_SIGNED(-25,11),
TO_SIGNED(-71,11),
TO_SIGNED(-118,11),
TO_SIGNED(-164,11),
TO_SIGNED(-210,11),
TO_SIGNED(-255,11),
TO_SIGNED(-298,11),
TO_SIGNED(-341,11),
TO_SIGNED(-382,11),
TO_SIGNED(-422,11),
TO_SIGNED(-460,11),
TO_SIGNED(-496,11),
TO_SIGNED(-530,11),
TO_SIGNED(-562,11),
TO_SIGNED(-592,11),
TO_SIGNED(-620,11),
TO_SIGNED(-645,11),
TO_SIGNED(-668,11),
TO_SIGNED(-688,11),
TO_SIGNED(-705,11),
TO_SIGNED(-720,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-721,11),
TO_SIGNED(-706,11),
TO_SIGNED(-689,11),
TO_SIGNED(-669,11),
TO_SIGNED(-647,11),
TO_SIGNED(-622,11),
TO_SIGNED(-594,11),
TO_SIGNED(-564,11),
TO_SIGNED(-532,11),
TO_SIGNED(-498,11),
TO_SIGNED(-462,11),
TO_SIGNED(-424,11),
TO_SIGNED(-385,11),
TO_SIGNED(-344,11),
TO_SIGNED(-301,11),
TO_SIGNED(-258,11),
TO_SIGNED(-213,11),
TO_SIGNED(-167,11),
TO_SIGNED(-121,11),
TO_SIGNED(-75,11),
TO_SIGNED(-28,11),
TO_SIGNED(19,11),
TO_SIGNED(66,11),
TO_SIGNED(113,11),
TO_SIGNED(159,11),
TO_SIGNED(205,11),
TO_SIGNED(249,11),
TO_SIGNED(293,11),
TO_SIGNED(336,11),
TO_SIGNED(377,11),
TO_SIGNED(417,11),
TO_SIGNED(455,11),
TO_SIGNED(492,11),
TO_SIGNED(526,11),
TO_SIGNED(559,11),
TO_SIGNED(589,11),
TO_SIGNED(617,11),
TO_SIGNED(642,11),
TO_SIGNED(665,11),
TO_SIGNED(686,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(708,11),
TO_SIGNED(691,11),
TO_SIGNED(672,11),
TO_SIGNED(650,11),
TO_SIGNED(625,11),
TO_SIGNED(598,11),
TO_SIGNED(568,11),
TO_SIGNED(536,11),
TO_SIGNED(502,11),
TO_SIGNED(466,11),
TO_SIGNED(429,11),
TO_SIGNED(389,11),
TO_SIGNED(348,11),
TO_SIGNED(306,11),
TO_SIGNED(263,11),
TO_SIGNED(218,11),
TO_SIGNED(173,11),
TO_SIGNED(127,11),
TO_SIGNED(80,11),
TO_SIGNED(33,11),
TO_SIGNED(-14,11),
TO_SIGNED(-61,11),
TO_SIGNED(-108,11),
TO_SIGNED(-154,11),
TO_SIGNED(-200,11),
TO_SIGNED(-244,11),
TO_SIGNED(-288,11),
TO_SIGNED(-331,11),
TO_SIGNED(-373,11),
TO_SIGNED(-413,11),
TO_SIGNED(-451,11),
TO_SIGNED(-488,11),
TO_SIGNED(-523,11),
TO_SIGNED(-555,11),
TO_SIGNED(-586,11),
TO_SIGNED(-614,11),
TO_SIGNED(-640,11),
TO_SIGNED(-663,11),
TO_SIGNED(-684,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-729,11),
TO_SIGNED(-739,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-710,11),
TO_SIGNED(-693,11),
TO_SIGNED(-674,11),
TO_SIGNED(-652,11),
TO_SIGNED(-628,11),
TO_SIGNED(-601,11),
TO_SIGNED(-571,11),
TO_SIGNED(-540,11),
TO_SIGNED(-506,11),
TO_SIGNED(-471,11),
TO_SIGNED(-433,11),
TO_SIGNED(-394,11),
TO_SIGNED(-353,11),
TO_SIGNED(-311,11),
TO_SIGNED(-268,11),
TO_SIGNED(-223,11),
TO_SIGNED(-178,11),
TO_SIGNED(-132,11),
TO_SIGNED(-85,11),
TO_SIGNED(-38,11),
TO_SIGNED(9,11),
TO_SIGNED(56,11),
TO_SIGNED(102,11),
TO_SIGNED(149,11),
TO_SIGNED(194,11),
TO_SIGNED(239,11),
TO_SIGNED(283,11),
TO_SIGNED(326,11),
TO_SIGNED(368,11),
TO_SIGNED(408,11),
TO_SIGNED(447,11),
TO_SIGNED(484,11),
TO_SIGNED(519,11),
TO_SIGNED(552,11),
TO_SIGNED(582,11),
TO_SIGNED(611,11),
TO_SIGNED(637,11),
TO_SIGNED(660,11),
TO_SIGNED(681,11),
TO_SIGNED(700,11),
TO_SIGNED(715,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(736,11),
TO_SIGNED(725,11),
TO_SIGNED(712,11),
TO_SIGNED(695,11),
TO_SIGNED(676,11),
TO_SIGNED(655,11),
TO_SIGNED(631,11),
TO_SIGNED(604,11),
TO_SIGNED(575,11),
TO_SIGNED(544,11),
TO_SIGNED(510,11),
TO_SIGNED(475,11),
TO_SIGNED(437,11),
TO_SIGNED(398,11),
TO_SIGNED(358,11),
TO_SIGNED(316,11),
TO_SIGNED(273,11),
TO_SIGNED(228,11),
TO_SIGNED(183,11),
TO_SIGNED(137,11),
TO_SIGNED(91,11),
TO_SIGNED(44,11),
TO_SIGNED(-3,11),
TO_SIGNED(-50,11),
TO_SIGNED(-97,11),
TO_SIGNED(-143,11),
TO_SIGNED(-189,11),
TO_SIGNED(-234,11),
TO_SIGNED(-278,11),
TO_SIGNED(-322,11),
TO_SIGNED(-363,11),
TO_SIGNED(-404,11),
TO_SIGNED(-443,11),
TO_SIGNED(-480,11),
TO_SIGNED(-515,11),
TO_SIGNED(-548,11),
TO_SIGNED(-579,11),
TO_SIGNED(-608,11),
TO_SIGNED(-634,11),
TO_SIGNED(-658,11),
TO_SIGNED(-679,11),
TO_SIGNED(-698,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-679,11),
TO_SIGNED(-657,11),
TO_SIGNED(-633,11),
TO_SIGNED(-607,11),
TO_SIGNED(-578,11),
TO_SIGNED(-547,11),
TO_SIGNED(-514,11),
TO_SIGNED(-479,11),
TO_SIGNED(-442,11),
TO_SIGNED(-403,11),
TO_SIGNED(-362,11),
TO_SIGNED(-321,11),
TO_SIGNED(-277,11),
TO_SIGNED(-233,11),
TO_SIGNED(-188,11),
TO_SIGNED(-142,11),
TO_SIGNED(-96,11),
TO_SIGNED(-49,11),
TO_SIGNED(-2,11),
TO_SIGNED(45,11),
TO_SIGNED(92,11),
TO_SIGNED(138,11),
TO_SIGNED(184,11),
TO_SIGNED(229,11),
TO_SIGNED(274,11),
TO_SIGNED(317,11),
TO_SIGNED(359,11),
TO_SIGNED(399,11),
TO_SIGNED(438,11),
TO_SIGNED(476,11),
TO_SIGNED(511,11),
TO_SIGNED(544,11),
TO_SIGNED(576,11),
TO_SIGNED(605,11),
TO_SIGNED(631,11),
TO_SIGNED(655,11),
TO_SIGNED(677,11),
TO_SIGNED(696,11),
TO_SIGNED(712,11),
TO_SIGNED(725,11),
TO_SIGNED(736,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(715,11),
TO_SIGNED(699,11),
TO_SIGNED(681,11),
TO_SIGNED(660,11),
TO_SIGNED(636,11),
TO_SIGNED(610,11),
TO_SIGNED(582,11),
TO_SIGNED(551,11),
TO_SIGNED(518,11),
TO_SIGNED(483,11),
TO_SIGNED(446,11),
TO_SIGNED(407,11),
TO_SIGNED(367,11),
TO_SIGNED(325,11),
TO_SIGNED(282,11),
TO_SIGNED(238,11),
TO_SIGNED(193,11),
TO_SIGNED(148,11),
TO_SIGNED(101,11),
TO_SIGNED(54,11),
TO_SIGNED(7,11),
TO_SIGNED(-40,11),
TO_SIGNED(-86,11),
TO_SIGNED(-133,11),
TO_SIGNED(-179,11),
TO_SIGNED(-224,11),
TO_SIGNED(-269,11),
TO_SIGNED(-312,11),
TO_SIGNED(-354,11),
TO_SIGNED(-395,11),
TO_SIGNED(-434,11),
TO_SIGNED(-471,11),
TO_SIGNED(-507,11),
TO_SIGNED(-541,11),
TO_SIGNED(-572,11),
TO_SIGNED(-601,11),
TO_SIGNED(-628,11),
TO_SIGNED(-653,11),
TO_SIGNED(-675,11),
TO_SIGNED(-694,11),
TO_SIGNED(-710,11),
TO_SIGNED(-724,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-701,11),
TO_SIGNED(-683,11),
TO_SIGNED(-662,11),
TO_SIGNED(-639,11),
TO_SIGNED(-613,11),
TO_SIGNED(-585,11),
TO_SIGNED(-554,11),
TO_SIGNED(-522,11),
TO_SIGNED(-487,11),
TO_SIGNED(-450,11),
TO_SIGNED(-412,11),
TO_SIGNED(-372,11),
TO_SIGNED(-330,11),
TO_SIGNED(-287,11),
TO_SIGNED(-243,11),
TO_SIGNED(-198,11),
TO_SIGNED(-153,11),
TO_SIGNED(-106,11),
TO_SIGNED(-60,11),
TO_SIGNED(-13,11),
TO_SIGNED(34,11),
TO_SIGNED(81,11),
TO_SIGNED(128,11),
TO_SIGNED(174,11),
TO_SIGNED(219,11),
TO_SIGNED(264,11),
TO_SIGNED(307,11),
TO_SIGNED(349,11),
TO_SIGNED(390,11),
TO_SIGNED(430,11),
TO_SIGNED(467,11),
TO_SIGNED(503,11),
TO_SIGNED(537,11),
TO_SIGNED(569,11),
TO_SIGNED(598,11),
TO_SIGNED(625,11),
TO_SIGNED(650,11),
TO_SIGNED(672,11),
TO_SIGNED(692,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(730,11),
TO_SIGNED(718,11),
TO_SIGNED(703,11),
TO_SIGNED(685,11),
TO_SIGNED(665,11),
TO_SIGNED(642,11),
TO_SIGNED(616,11),
TO_SIGNED(588,11),
TO_SIGNED(558,11),
TO_SIGNED(526,11),
TO_SIGNED(491,11),
TO_SIGNED(455,11),
TO_SIGNED(416,11),
TO_SIGNED(376,11),
TO_SIGNED(335,11),
TO_SIGNED(292,11),
TO_SIGNED(248,11),
TO_SIGNED(204,11),
TO_SIGNED(158,11),
TO_SIGNED(112,11),
TO_SIGNED(65,11),
TO_SIGNED(18,11),
TO_SIGNED(-29,11),
TO_SIGNED(-76,11),
TO_SIGNED(-122,11),
TO_SIGNED(-168,11),
TO_SIGNED(-214,11),
TO_SIGNED(-259,11),
TO_SIGNED(-302,11),
TO_SIGNED(-345,11),
TO_SIGNED(-386,11),
TO_SIGNED(-425,11),
TO_SIGNED(-463,11),
TO_SIGNED(-499,11),
TO_SIGNED(-533,11),
TO_SIGNED(-565,11),
TO_SIGNED(-595,11),
TO_SIGNED(-622,11),
TO_SIGNED(-647,11),
TO_SIGNED(-670,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-721,11),
TO_SIGNED(-733,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-720,11),
TO_SIGNED(-705,11),
TO_SIGNED(-688,11),
TO_SIGNED(-667,11),
TO_SIGNED(-645,11),
TO_SIGNED(-619,11),
TO_SIGNED(-592,11),
TO_SIGNED(-562,11),
TO_SIGNED(-529,11),
TO_SIGNED(-495,11),
TO_SIGNED(-459,11),
TO_SIGNED(-421,11),
TO_SIGNED(-381,11),
TO_SIGNED(-340,11),
TO_SIGNED(-297,11),
TO_SIGNED(-254,11),
TO_SIGNED(-209,11),
TO_SIGNED(-163,11),
TO_SIGNED(-117,11),
TO_SIGNED(-70,11),
TO_SIGNED(-24,11),
TO_SIGNED(24,11),
TO_SIGNED(70,11),
TO_SIGNED(117,11),
TO_SIGNED(163,11),
TO_SIGNED(209,11),
TO_SIGNED(254,11),
TO_SIGNED(297,11),
TO_SIGNED(340,11),
TO_SIGNED(381,11),
TO_SIGNED(421,11),
TO_SIGNED(459,11),
TO_SIGNED(495,11),
TO_SIGNED(529,11),
TO_SIGNED(562,11),
TO_SIGNED(592,11),
TO_SIGNED(619,11),
TO_SIGNED(645,11),
TO_SIGNED(667,11),
TO_SIGNED(688,11),
TO_SIGNED(705,11),
TO_SIGNED(720,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(733,11),
TO_SIGNED(721,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(670,11),
TO_SIGNED(647,11),
TO_SIGNED(622,11),
TO_SIGNED(595,11),
TO_SIGNED(565,11),
TO_SIGNED(533,11),
TO_SIGNED(499,11),
TO_SIGNED(463,11),
TO_SIGNED(425,11),
TO_SIGNED(386,11),
TO_SIGNED(345,11),
TO_SIGNED(302,11),
TO_SIGNED(259,11),
TO_SIGNED(214,11),
TO_SIGNED(168,11),
TO_SIGNED(122,11),
TO_SIGNED(76,11),
TO_SIGNED(29,11),
TO_SIGNED(-18,11),
TO_SIGNED(-65,11),
TO_SIGNED(-112,11),
TO_SIGNED(-158,11),
TO_SIGNED(-204,11),
TO_SIGNED(-248,11),
TO_SIGNED(-292,11),
TO_SIGNED(-335,11),
TO_SIGNED(-376,11),
TO_SIGNED(-416,11),
TO_SIGNED(-455,11),
TO_SIGNED(-491,11),
TO_SIGNED(-526,11),
TO_SIGNED(-558,11),
TO_SIGNED(-588,11),
TO_SIGNED(-616,11),
TO_SIGNED(-642,11),
TO_SIGNED(-665,11),
TO_SIGNED(-685,11),
TO_SIGNED(-703,11),
TO_SIGNED(-718,11),
TO_SIGNED(-730,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-692,11),
TO_SIGNED(-672,11),
TO_SIGNED(-650,11),
TO_SIGNED(-625,11),
TO_SIGNED(-598,11),
TO_SIGNED(-569,11),
TO_SIGNED(-537,11),
TO_SIGNED(-503,11),
TO_SIGNED(-467,11),
TO_SIGNED(-430,11),
TO_SIGNED(-390,11),
TO_SIGNED(-349,11),
TO_SIGNED(-307,11),
TO_SIGNED(-264,11),
TO_SIGNED(-219,11),
TO_SIGNED(-174,11),
TO_SIGNED(-128,11),
TO_SIGNED(-81,11),
TO_SIGNED(-34,11),
TO_SIGNED(13,11),
TO_SIGNED(60,11),
TO_SIGNED(106,11),
TO_SIGNED(153,11),
TO_SIGNED(198,11),
TO_SIGNED(243,11),
TO_SIGNED(287,11),
TO_SIGNED(330,11),
TO_SIGNED(372,11),
TO_SIGNED(412,11),
TO_SIGNED(450,11),
TO_SIGNED(487,11),
TO_SIGNED(522,11),
TO_SIGNED(554,11),
TO_SIGNED(585,11),
TO_SIGNED(613,11),
TO_SIGNED(639,11),
TO_SIGNED(662,11),
TO_SIGNED(683,11),
TO_SIGNED(701,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(724,11),
TO_SIGNED(710,11),
TO_SIGNED(694,11),
TO_SIGNED(675,11),
TO_SIGNED(653,11),
TO_SIGNED(628,11),
TO_SIGNED(601,11),
TO_SIGNED(572,11),
TO_SIGNED(541,11),
TO_SIGNED(507,11),
TO_SIGNED(471,11),
TO_SIGNED(434,11),
TO_SIGNED(395,11),
TO_SIGNED(354,11),
TO_SIGNED(312,11),
TO_SIGNED(269,11),
TO_SIGNED(224,11),
TO_SIGNED(179,11),
TO_SIGNED(133,11),
TO_SIGNED(86,11),
TO_SIGNED(40,11),
TO_SIGNED(-7,11),
TO_SIGNED(-54,11),
TO_SIGNED(-101,11),
TO_SIGNED(-148,11),
TO_SIGNED(-193,11),
TO_SIGNED(-238,11),
TO_SIGNED(-282,11),
TO_SIGNED(-325,11),
TO_SIGNED(-367,11),
TO_SIGNED(-407,11),
TO_SIGNED(-446,11),
TO_SIGNED(-483,11),
TO_SIGNED(-518,11),
TO_SIGNED(-551,11),
TO_SIGNED(-582,11),
TO_SIGNED(-610,11),
TO_SIGNED(-636,11),
TO_SIGNED(-660,11),
TO_SIGNED(-681,11),
TO_SIGNED(-699,11),
TO_SIGNED(-715,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-736,11),
TO_SIGNED(-725,11),
TO_SIGNED(-712,11),
TO_SIGNED(-696,11),
TO_SIGNED(-677,11),
TO_SIGNED(-655,11),
TO_SIGNED(-631,11),
TO_SIGNED(-605,11),
TO_SIGNED(-576,11),
TO_SIGNED(-544,11),
TO_SIGNED(-511,11),
TO_SIGNED(-476,11),
TO_SIGNED(-438,11),
TO_SIGNED(-399,11),
TO_SIGNED(-359,11),
TO_SIGNED(-317,11),
TO_SIGNED(-274,11),
TO_SIGNED(-229,11),
TO_SIGNED(-184,11),
TO_SIGNED(-138,11),
TO_SIGNED(-92,11),
TO_SIGNED(-45,11),
TO_SIGNED(2,11),
TO_SIGNED(49,11),
TO_SIGNED(96,11),
TO_SIGNED(142,11),
TO_SIGNED(188,11),
TO_SIGNED(233,11),
TO_SIGNED(277,11),
TO_SIGNED(321,11),
TO_SIGNED(362,11),
TO_SIGNED(403,11),
TO_SIGNED(442,11),
TO_SIGNED(479,11),
TO_SIGNED(514,11),
TO_SIGNED(547,11),
TO_SIGNED(578,11),
TO_SIGNED(607,11),
TO_SIGNED(633,11),
TO_SIGNED(657,11),
TO_SIGNED(679,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(698,11),
TO_SIGNED(679,11),
TO_SIGNED(658,11),
TO_SIGNED(634,11),
TO_SIGNED(608,11),
TO_SIGNED(579,11),
TO_SIGNED(548,11),
TO_SIGNED(515,11),
TO_SIGNED(480,11),
TO_SIGNED(443,11),
TO_SIGNED(404,11),
TO_SIGNED(363,11),
TO_SIGNED(322,11),
TO_SIGNED(278,11),
TO_SIGNED(234,11),
TO_SIGNED(189,11),
TO_SIGNED(143,11),
TO_SIGNED(97,11),
TO_SIGNED(50,11),
TO_SIGNED(3,11),
TO_SIGNED(-44,11),
TO_SIGNED(-91,11),
TO_SIGNED(-137,11),
TO_SIGNED(-183,11),
TO_SIGNED(-228,11),
TO_SIGNED(-273,11),
TO_SIGNED(-316,11),
TO_SIGNED(-358,11),
TO_SIGNED(-398,11),
TO_SIGNED(-437,11),
TO_SIGNED(-475,11),
TO_SIGNED(-510,11),
TO_SIGNED(-544,11),
TO_SIGNED(-575,11),
TO_SIGNED(-604,11),
TO_SIGNED(-631,11),
TO_SIGNED(-655,11),
TO_SIGNED(-676,11),
TO_SIGNED(-695,11),
TO_SIGNED(-712,11),
TO_SIGNED(-725,11),
TO_SIGNED(-736,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-715,11),
TO_SIGNED(-700,11),
TO_SIGNED(-681,11),
TO_SIGNED(-660,11),
TO_SIGNED(-637,11),
TO_SIGNED(-611,11),
TO_SIGNED(-582,11),
TO_SIGNED(-552,11),
TO_SIGNED(-519,11),
TO_SIGNED(-484,11),
TO_SIGNED(-447,11),
TO_SIGNED(-408,11),
TO_SIGNED(-368,11),
TO_SIGNED(-326,11),
TO_SIGNED(-283,11),
TO_SIGNED(-239,11),
TO_SIGNED(-194,11),
TO_SIGNED(-149,11),
TO_SIGNED(-102,11),
TO_SIGNED(-56,11),
TO_SIGNED(-9,11),
TO_SIGNED(38,11),
TO_SIGNED(85,11),
TO_SIGNED(132,11),
TO_SIGNED(178,11),
TO_SIGNED(223,11),
TO_SIGNED(268,11),
TO_SIGNED(311,11),
TO_SIGNED(353,11),
TO_SIGNED(394,11),
TO_SIGNED(433,11),
TO_SIGNED(471,11),
TO_SIGNED(506,11),
TO_SIGNED(540,11),
TO_SIGNED(571,11),
TO_SIGNED(601,11),
TO_SIGNED(628,11),
TO_SIGNED(652,11),
TO_SIGNED(674,11),
TO_SIGNED(693,11),
TO_SIGNED(710,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(739,11),
TO_SIGNED(729,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(684,11),
TO_SIGNED(663,11),
TO_SIGNED(640,11),
TO_SIGNED(614,11),
TO_SIGNED(586,11),
TO_SIGNED(555,11),
TO_SIGNED(523,11),
TO_SIGNED(488,11),
TO_SIGNED(451,11),
TO_SIGNED(413,11),
TO_SIGNED(373,11),
TO_SIGNED(331,11),
TO_SIGNED(288,11),
TO_SIGNED(244,11),
TO_SIGNED(200,11),
TO_SIGNED(154,11),
TO_SIGNED(108,11),
TO_SIGNED(61,11),
TO_SIGNED(14,11),
TO_SIGNED(-33,11),
TO_SIGNED(-80,11),
TO_SIGNED(-127,11),
TO_SIGNED(-173,11),
TO_SIGNED(-218,11),
TO_SIGNED(-263,11),
TO_SIGNED(-306,11),
TO_SIGNED(-348,11),
TO_SIGNED(-389,11),
TO_SIGNED(-429,11),
TO_SIGNED(-466,11),
TO_SIGNED(-502,11),
TO_SIGNED(-536,11),
TO_SIGNED(-568,11),
TO_SIGNED(-598,11),
TO_SIGNED(-625,11),
TO_SIGNED(-650,11),
TO_SIGNED(-672,11),
TO_SIGNED(-691,11),
TO_SIGNED(-708,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-686,11),
TO_SIGNED(-665,11),
TO_SIGNED(-642,11),
TO_SIGNED(-617,11),
TO_SIGNED(-589,11),
TO_SIGNED(-559,11),
TO_SIGNED(-526,11),
TO_SIGNED(-492,11),
TO_SIGNED(-455,11),
TO_SIGNED(-417,11),
TO_SIGNED(-377,11),
TO_SIGNED(-336,11),
TO_SIGNED(-293,11),
TO_SIGNED(-249,11),
TO_SIGNED(-205,11),
TO_SIGNED(-159,11),
TO_SIGNED(-113,11),
TO_SIGNED(-66,11),
TO_SIGNED(-19,11),
TO_SIGNED(28,11),
TO_SIGNED(75,11),
TO_SIGNED(121,11),
TO_SIGNED(167,11),
TO_SIGNED(213,11),
TO_SIGNED(258,11),
TO_SIGNED(301,11),
TO_SIGNED(344,11),
TO_SIGNED(385,11),
TO_SIGNED(424,11),
TO_SIGNED(462,11),
TO_SIGNED(498,11),
TO_SIGNED(532,11),
TO_SIGNED(564,11),
TO_SIGNED(594,11),
TO_SIGNED(622,11),
TO_SIGNED(647,11),
TO_SIGNED(669,11),
TO_SIGNED(689,11),
TO_SIGNED(706,11),
TO_SIGNED(721,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(720,11),
TO_SIGNED(705,11),
TO_SIGNED(688,11),
TO_SIGNED(668,11),
TO_SIGNED(645,11),
TO_SIGNED(620,11),
TO_SIGNED(592,11),
TO_SIGNED(562,11),
TO_SIGNED(530,11),
TO_SIGNED(496,11),
TO_SIGNED(460,11),
TO_SIGNED(422,11),
TO_SIGNED(382,11),
TO_SIGNED(341,11),
TO_SIGNED(298,11),
TO_SIGNED(255,11),
TO_SIGNED(210,11),
TO_SIGNED(164,11),
TO_SIGNED(118,11),
TO_SIGNED(71,11),
TO_SIGNED(25,11),
TO_SIGNED(-22,11),
TO_SIGNED(-69,11),
TO_SIGNED(-116,11),
TO_SIGNED(-162,11),
TO_SIGNED(-208,11),
TO_SIGNED(-252,11),
TO_SIGNED(-296,11),
TO_SIGNED(-339,11),
TO_SIGNED(-380,11),
TO_SIGNED(-420,11),
TO_SIGNED(-458,11),
TO_SIGNED(-494,11),
TO_SIGNED(-529,11),
TO_SIGNED(-561,11),
TO_SIGNED(-591,11),
TO_SIGNED(-619,11),
TO_SIGNED(-644,11),
TO_SIGNED(-667,11),
TO_SIGNED(-687,11),
TO_SIGNED(-705,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-733,11),
TO_SIGNED(-721,11),
TO_SIGNED(-707,11),
TO_SIGNED(-690,11),
TO_SIGNED(-670,11),
TO_SIGNED(-648,11),
TO_SIGNED(-623,11),
TO_SIGNED(-596,11),
TO_SIGNED(-566,11),
TO_SIGNED(-534,11),
TO_SIGNED(-500,11),
TO_SIGNED(-464,11),
TO_SIGNED(-426,11),
TO_SIGNED(-387,11),
TO_SIGNED(-345,11),
TO_SIGNED(-303,11),
TO_SIGNED(-260,11),
TO_SIGNED(-215,11),
TO_SIGNED(-169,11),
TO_SIGNED(-123,11),
TO_SIGNED(-77,11),
TO_SIGNED(-30,11),
TO_SIGNED(17,11),
TO_SIGNED(64,11),
TO_SIGNED(111,11),
TO_SIGNED(157,11),
TO_SIGNED(203,11),
TO_SIGNED(247,11),
TO_SIGNED(291,11),
TO_SIGNED(334,11),
TO_SIGNED(375,11),
TO_SIGNED(415,11),
TO_SIGNED(454,11),
TO_SIGNED(490,11),
TO_SIGNED(525,11),
TO_SIGNED(557,11),
TO_SIGNED(588,11),
TO_SIGNED(616,11),
TO_SIGNED(641,11),
TO_SIGNED(664,11),
TO_SIGNED(685,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(709,11),
TO_SIGNED(692,11),
TO_SIGNED(673,11),
TO_SIGNED(651,11),
TO_SIGNED(626,11),
TO_SIGNED(599,11),
TO_SIGNED(569,11),
TO_SIGNED(538,11),
TO_SIGNED(504,11),
TO_SIGNED(468,11),
TO_SIGNED(430,11),
TO_SIGNED(391,11),
TO_SIGNED(350,11),
TO_SIGNED(308,11),
TO_SIGNED(265,11),
TO_SIGNED(220,11),
TO_SIGNED(175,11),
TO_SIGNED(129,11),
TO_SIGNED(82,11),
TO_SIGNED(35,11),
TO_SIGNED(-12,11),
TO_SIGNED(-59,11),
TO_SIGNED(-105,11),
TO_SIGNED(-152,11),
TO_SIGNED(-197,11),
TO_SIGNED(-242,11),
TO_SIGNED(-286,11),
TO_SIGNED(-329,11),
TO_SIGNED(-371,11),
TO_SIGNED(-411,11),
TO_SIGNED(-449,11),
TO_SIGNED(-486,11),
TO_SIGNED(-521,11),
TO_SIGNED(-554,11),
TO_SIGNED(-584,11),
TO_SIGNED(-613,11),
TO_SIGNED(-639,11),
TO_SIGNED(-662,11),
TO_SIGNED(-683,11),
TO_SIGNED(-701,11),
TO_SIGNED(-716,11),
TO_SIGNED(-729,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-711,11),
TO_SIGNED(-694,11),
TO_SIGNED(-675,11),
TO_SIGNED(-653,11),
TO_SIGNED(-629,11),
TO_SIGNED(-602,11),
TO_SIGNED(-573,11),
TO_SIGNED(-541,11),
TO_SIGNED(-508,11),
TO_SIGNED(-472,11),
TO_SIGNED(-435,11),
TO_SIGNED(-396,11),
TO_SIGNED(-355,11),
TO_SIGNED(-313,11),
TO_SIGNED(-270,11),
TO_SIGNED(-225,11),
TO_SIGNED(-180,11),
TO_SIGNED(-134,11),
TO_SIGNED(-87,11),
TO_SIGNED(-41,11),
TO_SIGNED(6,11),
TO_SIGNED(53,11),
TO_SIGNED(100,11),
TO_SIGNED(147,11),
TO_SIGNED(192,11),
TO_SIGNED(237,11),
TO_SIGNED(281,11),
TO_SIGNED(324,11),
TO_SIGNED(366,11),
TO_SIGNED(406,11),
TO_SIGNED(445,11),
TO_SIGNED(482,11),
TO_SIGNED(517,11),
TO_SIGNED(550,11),
TO_SIGNED(581,11),
TO_SIGNED(610,11),
TO_SIGNED(636,11),
TO_SIGNED(659,11),
TO_SIGNED(681,11),
TO_SIGNED(699,11),
TO_SIGNED(715,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(712,11),
TO_SIGNED(696,11),
TO_SIGNED(677,11),
TO_SIGNED(656,11),
TO_SIGNED(632,11),
TO_SIGNED(605,11),
TO_SIGNED(576,11),
TO_SIGNED(545,11),
TO_SIGNED(512,11),
TO_SIGNED(476,11),
TO_SIGNED(439,11),
TO_SIGNED(400,11),
TO_SIGNED(360,11),
TO_SIGNED(318,11),
TO_SIGNED(275,11),
TO_SIGNED(230,11),
TO_SIGNED(185,11),
TO_SIGNED(139,11),
TO_SIGNED(93,11),
TO_SIGNED(46,11),
TO_SIGNED(-1,11),
TO_SIGNED(-48,11),
TO_SIGNED(-95,11),
TO_SIGNED(-141,11),
TO_SIGNED(-187,11),
TO_SIGNED(-232,11),
TO_SIGNED(-276,11),
TO_SIGNED(-320,11),
TO_SIGNED(-362,11),
TO_SIGNED(-402,11),
TO_SIGNED(-441,11),
TO_SIGNED(-478,11),
TO_SIGNED(-513,11),
TO_SIGNED(-547,11),
TO_SIGNED(-578,11),
TO_SIGNED(-606,11),
TO_SIGNED(-633,11),
TO_SIGNED(-657,11),
TO_SIGNED(-678,11),
TO_SIGNED(-697,11),
TO_SIGNED(-713,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-714,11),
TO_SIGNED(-698,11),
TO_SIGNED(-680,11),
TO_SIGNED(-658,11),
TO_SIGNED(-635,11),
TO_SIGNED(-608,11),
TO_SIGNED(-580,11),
TO_SIGNED(-549,11),
TO_SIGNED(-516,11),
TO_SIGNED(-480,11),
TO_SIGNED(-443,11),
TO_SIGNED(-405,11),
TO_SIGNED(-364,11),
TO_SIGNED(-323,11),
TO_SIGNED(-279,11),
TO_SIGNED(-235,11),
TO_SIGNED(-190,11),
TO_SIGNED(-144,11),
TO_SIGNED(-98,11),
TO_SIGNED(-51,11),
TO_SIGNED(-4,11),
TO_SIGNED(43,11),
TO_SIGNED(90,11),
TO_SIGNED(136,11),
TO_SIGNED(182,11),
TO_SIGNED(227,11),
TO_SIGNED(272,11),
TO_SIGNED(315,11),
TO_SIGNED(357,11),
TO_SIGNED(397,11),
TO_SIGNED(437,11),
TO_SIGNED(474,11),
TO_SIGNED(509,11),
TO_SIGNED(543,11),
TO_SIGNED(574,11),
TO_SIGNED(603,11),
TO_SIGNED(630,11),
TO_SIGNED(654,11),
TO_SIGNED(676,11),
TO_SIGNED(695,11),
TO_SIGNED(711,11),
TO_SIGNED(725,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(716,11),
TO_SIGNED(700,11),
TO_SIGNED(682,11),
TO_SIGNED(661,11),
TO_SIGNED(637,11),
TO_SIGNED(611,11),
TO_SIGNED(583,11),
TO_SIGNED(552,11),
TO_SIGNED(519,11),
TO_SIGNED(485,11),
TO_SIGNED(448,11),
TO_SIGNED(409,11),
TO_SIGNED(369,11),
TO_SIGNED(327,11),
TO_SIGNED(284,11),
TO_SIGNED(240,11),
TO_SIGNED(195,11),
TO_SIGNED(150,11),
TO_SIGNED(103,11),
TO_SIGNED(57,11),
TO_SIGNED(10,11),
TO_SIGNED(-37,11),
TO_SIGNED(-84,11),
TO_SIGNED(-131,11),
TO_SIGNED(-177,11),
TO_SIGNED(-222,11),
TO_SIGNED(-267,11),
TO_SIGNED(-310,11),
TO_SIGNED(-352,11),
TO_SIGNED(-393,11),
TO_SIGNED(-432,11),
TO_SIGNED(-470,11),
TO_SIGNED(-505,11),
TO_SIGNED(-539,11),
TO_SIGNED(-571,11),
TO_SIGNED(-600,11),
TO_SIGNED(-627,11),
TO_SIGNED(-652,11),
TO_SIGNED(-674,11),
TO_SIGNED(-693,11),
TO_SIGNED(-710,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-702,11),
TO_SIGNED(-684,11),
TO_SIGNED(-663,11),
TO_SIGNED(-640,11),
TO_SIGNED(-615,11),
TO_SIGNED(-586,11),
TO_SIGNED(-556,11),
TO_SIGNED(-523,11),
TO_SIGNED(-489,11),
TO_SIGNED(-452,11),
TO_SIGNED(-414,11),
TO_SIGNED(-374,11),
TO_SIGNED(-332,11),
TO_SIGNED(-289,11),
TO_SIGNED(-245,11),
TO_SIGNED(-201,11),
TO_SIGNED(-155,11),
TO_SIGNED(-109,11),
TO_SIGNED(-62,11),
TO_SIGNED(-15,11),
TO_SIGNED(32,11),
TO_SIGNED(79,11),
TO_SIGNED(125,11),
TO_SIGNED(172,11),
TO_SIGNED(217,11),
TO_SIGNED(262,11),
TO_SIGNED(305,11),
TO_SIGNED(347,11),
TO_SIGNED(388,11),
TO_SIGNED(428,11),
TO_SIGNED(466,11),
TO_SIGNED(501,11),
TO_SIGNED(535,11),
TO_SIGNED(567,11),
TO_SIGNED(597,11),
TO_SIGNED(624,11),
TO_SIGNED(649,11),
TO_SIGNED(671,11),
TO_SIGNED(691,11),
TO_SIGNED(708,11),
TO_SIGNED(722,11),
TO_SIGNED(733,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(704,11),
TO_SIGNED(686,11),
TO_SIGNED(666,11),
TO_SIGNED(643,11),
TO_SIGNED(618,11),
TO_SIGNED(590,11),
TO_SIGNED(559,11),
TO_SIGNED(527,11),
TO_SIGNED(493,11),
TO_SIGNED(456,11),
TO_SIGNED(418,11),
TO_SIGNED(378,11),
TO_SIGNED(337,11),
TO_SIGNED(294,11),
TO_SIGNED(250,11),
TO_SIGNED(206,11),
TO_SIGNED(160,11),
TO_SIGNED(114,11),
TO_SIGNED(67,11),
TO_SIGNED(20,11),
TO_SIGNED(-27,11),
TO_SIGNED(-74,11),
TO_SIGNED(-120,11),
TO_SIGNED(-166,11),
TO_SIGNED(-212,11),
TO_SIGNED(-257,11),
TO_SIGNED(-300,11),
TO_SIGNED(-343,11),
TO_SIGNED(-384,11),
TO_SIGNED(-423,11),
TO_SIGNED(-461,11),
TO_SIGNED(-497,11),
TO_SIGNED(-532,11),
TO_SIGNED(-564,11),
TO_SIGNED(-594,11),
TO_SIGNED(-621,11),
TO_SIGNED(-646,11),
TO_SIGNED(-669,11),
TO_SIGNED(-689,11),
TO_SIGNED(-706,11),
TO_SIGNED(-721,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-720,11),
TO_SIGNED(-706,11),
TO_SIGNED(-688,11),
TO_SIGNED(-668,11),
TO_SIGNED(-646,11),
TO_SIGNED(-621,11),
TO_SIGNED(-593,11),
TO_SIGNED(-563,11),
TO_SIGNED(-531,11),
TO_SIGNED(-497,11),
TO_SIGNED(-460,11),
TO_SIGNED(-422,11),
TO_SIGNED(-383,11),
TO_SIGNED(-342,11),
TO_SIGNED(-299,11),
TO_SIGNED(-256,11),
TO_SIGNED(-211,11),
TO_SIGNED(-165,11),
TO_SIGNED(-119,11),
TO_SIGNED(-73,11),
TO_SIGNED(-26,11),
TO_SIGNED(21,11),
TO_SIGNED(68,11),
TO_SIGNED(115,11),
TO_SIGNED(161,11),
TO_SIGNED(207,11),
TO_SIGNED(251,11),
TO_SIGNED(295,11),
TO_SIGNED(338,11),
TO_SIGNED(379,11),
TO_SIGNED(419,11),
TO_SIGNED(457,11),
TO_SIGNED(493,11),
TO_SIGNED(528,11),
TO_SIGNED(560,11),
TO_SIGNED(590,11),
TO_SIGNED(618,11),
TO_SIGNED(644,11),
TO_SIGNED(666,11),
TO_SIGNED(687,11),
TO_SIGNED(704,11),
TO_SIGNED(719,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(671,11),
TO_SIGNED(648,11),
TO_SIGNED(624,11),
TO_SIGNED(596,11),
TO_SIGNED(567,11),
TO_SIGNED(535,11),
TO_SIGNED(501,11),
TO_SIGNED(465,11),
TO_SIGNED(427,11),
TO_SIGNED(387,11),
TO_SIGNED(346,11),
TO_SIGNED(304,11),
TO_SIGNED(261,11),
TO_SIGNED(216,11),
TO_SIGNED(171,11),
TO_SIGNED(124,11),
TO_SIGNED(78,11),
TO_SIGNED(31,11),
TO_SIGNED(-16,11),
TO_SIGNED(-63,11),
TO_SIGNED(-110,11),
TO_SIGNED(-156,11),
TO_SIGNED(-202,11),
TO_SIGNED(-246,11),
TO_SIGNED(-290,11),
TO_SIGNED(-333,11),
TO_SIGNED(-375,11),
TO_SIGNED(-415,11),
TO_SIGNED(-453,11),
TO_SIGNED(-489,11),
TO_SIGNED(-524,11),
TO_SIGNED(-557,11),
TO_SIGNED(-587,11),
TO_SIGNED(-615,11),
TO_SIGNED(-641,11),
TO_SIGNED(-664,11),
TO_SIGNED(-685,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-730,11),
TO_SIGNED(-739,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-693,11),
TO_SIGNED(-673,11),
TO_SIGNED(-651,11),
TO_SIGNED(-627,11),
TO_SIGNED(-599,11),
TO_SIGNED(-570,11),
TO_SIGNED(-538,11),
TO_SIGNED(-505,11),
TO_SIGNED(-469,11),
TO_SIGNED(-431,11),
TO_SIGNED(-392,11),
TO_SIGNED(-351,11),
TO_SIGNED(-309,11),
TO_SIGNED(-266,11),
TO_SIGNED(-221,11),
TO_SIGNED(-176,11),
TO_SIGNED(-130,11),
TO_SIGNED(-83,11),
TO_SIGNED(-36,11),
TO_SIGNED(11,11),
TO_SIGNED(58,11),
TO_SIGNED(104,11),
TO_SIGNED(151,11),
TO_SIGNED(196,11),
TO_SIGNED(241,11),
TO_SIGNED(285,11),
TO_SIGNED(328,11),
TO_SIGNED(370,11),
TO_SIGNED(410,11),
TO_SIGNED(449,11),
TO_SIGNED(485,11),
TO_SIGNED(520,11),
TO_SIGNED(553,11),
TO_SIGNED(584,11),
TO_SIGNED(612,11),
TO_SIGNED(638,11),
TO_SIGNED(661,11),
TO_SIGNED(682,11),
TO_SIGNED(700,11),
TO_SIGNED(716,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(725,11),
TO_SIGNED(711,11),
TO_SIGNED(695,11),
TO_SIGNED(675,11),
TO_SIGNED(654,11),
TO_SIGNED(629,11),
TO_SIGNED(603,11),
TO_SIGNED(574,11),
TO_SIGNED(542,11),
TO_SIGNED(509,11),
TO_SIGNED(473,11),
TO_SIGNED(436,11),
TO_SIGNED(397,11),
TO_SIGNED(356,11),
TO_SIGNED(314,11),
TO_SIGNED(271,11),
TO_SIGNED(226,11),
TO_SIGNED(181,11),
TO_SIGNED(135,11),
TO_SIGNED(88,11),
TO_SIGNED(42,11),
TO_SIGNED(-5,11),
TO_SIGNED(-52,11),
TO_SIGNED(-99,11),
TO_SIGNED(-145,11),
TO_SIGNED(-191,11),
TO_SIGNED(-236,11),
TO_SIGNED(-280,11),
TO_SIGNED(-323,11),
TO_SIGNED(-365,11),
TO_SIGNED(-406,11),
TO_SIGNED(-444,11),
TO_SIGNED(-481,11),
TO_SIGNED(-516,11),
TO_SIGNED(-549,11),
TO_SIGNED(-580,11),
TO_SIGNED(-609,11),
TO_SIGNED(-635,11),
TO_SIGNED(-659,11),
TO_SIGNED(-680,11),
TO_SIGNED(-699,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-736,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-678,11),
TO_SIGNED(-656,11),
TO_SIGNED(-632,11),
TO_SIGNED(-606,11),
TO_SIGNED(-577,11),
TO_SIGNED(-546,11),
TO_SIGNED(-512,11),
TO_SIGNED(-477,11),
TO_SIGNED(-440,11),
TO_SIGNED(-401,11),
TO_SIGNED(-361,11),
TO_SIGNED(-319,11),
TO_SIGNED(-275,11),
TO_SIGNED(-231,11),
TO_SIGNED(-186,11),
TO_SIGNED(-140,11),
TO_SIGNED(-94,11),
TO_SIGNED(-47,11),
TO_SIGNED(0,11),
TO_SIGNED(47,11),
TO_SIGNED(94,11),
TO_SIGNED(140,11),
TO_SIGNED(186,11),
TO_SIGNED(231,11),
TO_SIGNED(275,11),
TO_SIGNED(319,11),
TO_SIGNED(361,11),
TO_SIGNED(401,11),
TO_SIGNED(440,11),
TO_SIGNED(477,11),
TO_SIGNED(512,11),
TO_SIGNED(546,11),
TO_SIGNED(577,11),
TO_SIGNED(606,11),
TO_SIGNED(632,11),
TO_SIGNED(656,11),
TO_SIGNED(678,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(736,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(699,11),
TO_SIGNED(680,11),
TO_SIGNED(659,11),
TO_SIGNED(635,11),
TO_SIGNED(609,11),
TO_SIGNED(580,11),
TO_SIGNED(549,11),
TO_SIGNED(516,11),
TO_SIGNED(481,11),
TO_SIGNED(444,11),
TO_SIGNED(406,11),
TO_SIGNED(365,11),
TO_SIGNED(323,11),
TO_SIGNED(280,11),
TO_SIGNED(236,11),
TO_SIGNED(191,11),
TO_SIGNED(145,11),
TO_SIGNED(99,11),
TO_SIGNED(52,11),
TO_SIGNED(5,11),
TO_SIGNED(-42,11),
TO_SIGNED(-88,11),
TO_SIGNED(-135,11),
TO_SIGNED(-181,11),
TO_SIGNED(-226,11),
TO_SIGNED(-271,11),
TO_SIGNED(-314,11),
TO_SIGNED(-356,11),
TO_SIGNED(-397,11),
TO_SIGNED(-436,11),
TO_SIGNED(-473,11),
TO_SIGNED(-509,11),
TO_SIGNED(-542,11),
TO_SIGNED(-574,11),
TO_SIGNED(-603,11),
TO_SIGNED(-629,11),
TO_SIGNED(-654,11),
TO_SIGNED(-675,11),
TO_SIGNED(-695,11),
TO_SIGNED(-711,11),
TO_SIGNED(-725,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-716,11),
TO_SIGNED(-700,11),
TO_SIGNED(-682,11),
TO_SIGNED(-661,11),
TO_SIGNED(-638,11),
TO_SIGNED(-612,11),
TO_SIGNED(-584,11),
TO_SIGNED(-553,11),
TO_SIGNED(-520,11),
TO_SIGNED(-485,11),
TO_SIGNED(-449,11),
TO_SIGNED(-410,11),
TO_SIGNED(-370,11),
TO_SIGNED(-328,11),
TO_SIGNED(-285,11),
TO_SIGNED(-241,11),
TO_SIGNED(-196,11),
TO_SIGNED(-151,11),
TO_SIGNED(-104,11),
TO_SIGNED(-58,11),
TO_SIGNED(-11,11),
TO_SIGNED(36,11),
TO_SIGNED(83,11),
TO_SIGNED(130,11),
TO_SIGNED(176,11),
TO_SIGNED(221,11),
TO_SIGNED(266,11),
TO_SIGNED(309,11),
TO_SIGNED(351,11),
TO_SIGNED(392,11),
TO_SIGNED(431,11),
TO_SIGNED(469,11),
TO_SIGNED(505,11),
TO_SIGNED(538,11),
TO_SIGNED(570,11),
TO_SIGNED(599,11),
TO_SIGNED(627,11),
TO_SIGNED(651,11),
TO_SIGNED(673,11),
TO_SIGNED(693,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(739,11),
TO_SIGNED(730,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(685,11),
TO_SIGNED(664,11),
TO_SIGNED(641,11),
TO_SIGNED(615,11),
TO_SIGNED(587,11),
TO_SIGNED(557,11),
TO_SIGNED(524,11),
TO_SIGNED(489,11),
TO_SIGNED(453,11),
TO_SIGNED(415,11),
TO_SIGNED(375,11),
TO_SIGNED(333,11),
TO_SIGNED(290,11),
TO_SIGNED(246,11),
TO_SIGNED(202,11),
TO_SIGNED(156,11),
TO_SIGNED(110,11),
TO_SIGNED(63,11),
TO_SIGNED(16,11),
TO_SIGNED(-31,11),
TO_SIGNED(-78,11),
TO_SIGNED(-124,11),
TO_SIGNED(-171,11),
TO_SIGNED(-216,11),
TO_SIGNED(-261,11),
TO_SIGNED(-304,11),
TO_SIGNED(-346,11),
TO_SIGNED(-387,11),
TO_SIGNED(-427,11),
TO_SIGNED(-465,11),
TO_SIGNED(-501,11),
TO_SIGNED(-535,11),
TO_SIGNED(-567,11),
TO_SIGNED(-596,11),
TO_SIGNED(-624,11),
TO_SIGNED(-648,11),
TO_SIGNED(-671,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-719,11),
TO_SIGNED(-704,11),
TO_SIGNED(-687,11),
TO_SIGNED(-666,11),
TO_SIGNED(-644,11),
TO_SIGNED(-618,11),
TO_SIGNED(-590,11),
TO_SIGNED(-560,11),
TO_SIGNED(-528,11),
TO_SIGNED(-493,11),
TO_SIGNED(-457,11),
TO_SIGNED(-419,11),
TO_SIGNED(-379,11),
TO_SIGNED(-338,11),
TO_SIGNED(-295,11),
TO_SIGNED(-251,11),
TO_SIGNED(-207,11),
TO_SIGNED(-161,11),
TO_SIGNED(-115,11),
TO_SIGNED(-68,11),
TO_SIGNED(-21,11),
TO_SIGNED(26,11),
TO_SIGNED(73,11),
TO_SIGNED(119,11),
TO_SIGNED(165,11),
TO_SIGNED(211,11),
TO_SIGNED(256,11),
TO_SIGNED(299,11),
TO_SIGNED(342,11),
TO_SIGNED(383,11),
TO_SIGNED(422,11),
TO_SIGNED(460,11),
TO_SIGNED(497,11),
TO_SIGNED(531,11),
TO_SIGNED(563,11),
TO_SIGNED(593,11),
TO_SIGNED(621,11),
TO_SIGNED(646,11),
TO_SIGNED(668,11),
TO_SIGNED(688,11),
TO_SIGNED(706,11),
TO_SIGNED(720,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(721,11),
TO_SIGNED(706,11),
TO_SIGNED(689,11),
TO_SIGNED(669,11),
TO_SIGNED(646,11),
TO_SIGNED(621,11),
TO_SIGNED(594,11),
TO_SIGNED(564,11),
TO_SIGNED(532,11),
TO_SIGNED(497,11),
TO_SIGNED(461,11),
TO_SIGNED(423,11),
TO_SIGNED(384,11),
TO_SIGNED(343,11),
TO_SIGNED(300,11),
TO_SIGNED(257,11),
TO_SIGNED(212,11),
TO_SIGNED(166,11),
TO_SIGNED(120,11),
TO_SIGNED(74,11),
TO_SIGNED(27,11),
TO_SIGNED(-20,11),
TO_SIGNED(-67,11),
TO_SIGNED(-114,11),
TO_SIGNED(-160,11),
TO_SIGNED(-206,11),
TO_SIGNED(-250,11),
TO_SIGNED(-294,11),
TO_SIGNED(-337,11),
TO_SIGNED(-378,11),
TO_SIGNED(-418,11),
TO_SIGNED(-456,11),
TO_SIGNED(-493,11),
TO_SIGNED(-527,11),
TO_SIGNED(-559,11),
TO_SIGNED(-590,11),
TO_SIGNED(-618,11),
TO_SIGNED(-643,11),
TO_SIGNED(-666,11),
TO_SIGNED(-686,11),
TO_SIGNED(-704,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-733,11),
TO_SIGNED(-722,11),
TO_SIGNED(-708,11),
TO_SIGNED(-691,11),
TO_SIGNED(-671,11),
TO_SIGNED(-649,11),
TO_SIGNED(-624,11),
TO_SIGNED(-597,11),
TO_SIGNED(-567,11),
TO_SIGNED(-535,11),
TO_SIGNED(-501,11),
TO_SIGNED(-466,11),
TO_SIGNED(-428,11),
TO_SIGNED(-388,11),
TO_SIGNED(-347,11),
TO_SIGNED(-305,11),
TO_SIGNED(-262,11),
TO_SIGNED(-217,11),
TO_SIGNED(-172,11),
TO_SIGNED(-125,11),
TO_SIGNED(-79,11),
TO_SIGNED(-32,11),
TO_SIGNED(15,11),
TO_SIGNED(62,11),
TO_SIGNED(109,11),
TO_SIGNED(155,11),
TO_SIGNED(201,11),
TO_SIGNED(245,11),
TO_SIGNED(289,11),
TO_SIGNED(332,11),
TO_SIGNED(374,11),
TO_SIGNED(414,11),
TO_SIGNED(452,11),
TO_SIGNED(489,11),
TO_SIGNED(523,11),
TO_SIGNED(556,11),
TO_SIGNED(586,11),
TO_SIGNED(615,11),
TO_SIGNED(640,11),
TO_SIGNED(663,11),
TO_SIGNED(684,11),
TO_SIGNED(702,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(710,11),
TO_SIGNED(693,11),
TO_SIGNED(674,11),
TO_SIGNED(652,11),
TO_SIGNED(627,11),
TO_SIGNED(600,11),
TO_SIGNED(571,11),
TO_SIGNED(539,11),
TO_SIGNED(505,11),
TO_SIGNED(470,11),
TO_SIGNED(432,11),
TO_SIGNED(393,11),
TO_SIGNED(352,11),
TO_SIGNED(310,11),
TO_SIGNED(267,11),
TO_SIGNED(222,11),
TO_SIGNED(177,11),
TO_SIGNED(131,11),
TO_SIGNED(84,11),
TO_SIGNED(37,11),
TO_SIGNED(-10,11),
TO_SIGNED(-57,11),
TO_SIGNED(-103,11),
TO_SIGNED(-150,11),
TO_SIGNED(-195,11),
TO_SIGNED(-240,11),
TO_SIGNED(-284,11),
TO_SIGNED(-327,11),
TO_SIGNED(-369,11),
TO_SIGNED(-409,11),
TO_SIGNED(-448,11),
TO_SIGNED(-485,11),
TO_SIGNED(-519,11),
TO_SIGNED(-552,11),
TO_SIGNED(-583,11),
TO_SIGNED(-611,11),
TO_SIGNED(-637,11),
TO_SIGNED(-661,11),
TO_SIGNED(-682,11),
TO_SIGNED(-700,11),
TO_SIGNED(-716,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-725,11),
TO_SIGNED(-711,11),
TO_SIGNED(-695,11),
TO_SIGNED(-676,11),
TO_SIGNED(-654,11),
TO_SIGNED(-630,11),
TO_SIGNED(-603,11),
TO_SIGNED(-574,11),
TO_SIGNED(-543,11),
TO_SIGNED(-509,11),
TO_SIGNED(-474,11),
TO_SIGNED(-437,11),
TO_SIGNED(-397,11),
TO_SIGNED(-357,11),
TO_SIGNED(-315,11),
TO_SIGNED(-272,11),
TO_SIGNED(-227,11),
TO_SIGNED(-182,11),
TO_SIGNED(-136,11),
TO_SIGNED(-90,11),
TO_SIGNED(-43,11),
TO_SIGNED(4,11),
TO_SIGNED(51,11),
TO_SIGNED(98,11),
TO_SIGNED(144,11),
TO_SIGNED(190,11),
TO_SIGNED(235,11),
TO_SIGNED(279,11),
TO_SIGNED(323,11),
TO_SIGNED(364,11),
TO_SIGNED(405,11),
TO_SIGNED(443,11),
TO_SIGNED(480,11),
TO_SIGNED(516,11),
TO_SIGNED(549,11),
TO_SIGNED(580,11),
TO_SIGNED(608,11),
TO_SIGNED(635,11),
TO_SIGNED(658,11),
TO_SIGNED(680,11),
TO_SIGNED(698,11),
TO_SIGNED(714,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(713,11),
TO_SIGNED(697,11),
TO_SIGNED(678,11),
TO_SIGNED(657,11),
TO_SIGNED(633,11),
TO_SIGNED(606,11),
TO_SIGNED(578,11),
TO_SIGNED(547,11),
TO_SIGNED(513,11),
TO_SIGNED(478,11),
TO_SIGNED(441,11),
TO_SIGNED(402,11),
TO_SIGNED(362,11),
TO_SIGNED(320,11),
TO_SIGNED(276,11),
TO_SIGNED(232,11),
TO_SIGNED(187,11),
TO_SIGNED(141,11),
TO_SIGNED(95,11),
TO_SIGNED(48,11),
TO_SIGNED(1,11),
TO_SIGNED(-46,11),
TO_SIGNED(-93,11),
TO_SIGNED(-139,11),
TO_SIGNED(-185,11),
TO_SIGNED(-230,11),
TO_SIGNED(-275,11),
TO_SIGNED(-318,11),
TO_SIGNED(-360,11),
TO_SIGNED(-400,11),
TO_SIGNED(-439,11),
TO_SIGNED(-476,11),
TO_SIGNED(-512,11),
TO_SIGNED(-545,11),
TO_SIGNED(-576,11),
TO_SIGNED(-605,11),
TO_SIGNED(-632,11),
TO_SIGNED(-656,11),
TO_SIGNED(-677,11),
TO_SIGNED(-696,11),
TO_SIGNED(-712,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-715,11),
TO_SIGNED(-699,11),
TO_SIGNED(-681,11),
TO_SIGNED(-659,11),
TO_SIGNED(-636,11),
TO_SIGNED(-610,11),
TO_SIGNED(-581,11),
TO_SIGNED(-550,11),
TO_SIGNED(-517,11),
TO_SIGNED(-482,11),
TO_SIGNED(-445,11),
TO_SIGNED(-406,11),
TO_SIGNED(-366,11),
TO_SIGNED(-324,11),
TO_SIGNED(-281,11),
TO_SIGNED(-237,11),
TO_SIGNED(-192,11),
TO_SIGNED(-147,11),
TO_SIGNED(-100,11),
TO_SIGNED(-53,11),
TO_SIGNED(-6,11),
TO_SIGNED(41,11),
TO_SIGNED(87,11),
TO_SIGNED(134,11),
TO_SIGNED(180,11),
TO_SIGNED(225,11),
TO_SIGNED(270,11),
TO_SIGNED(313,11),
TO_SIGNED(355,11),
TO_SIGNED(396,11),
TO_SIGNED(435,11),
TO_SIGNED(472,11),
TO_SIGNED(508,11),
TO_SIGNED(541,11),
TO_SIGNED(573,11),
TO_SIGNED(602,11),
TO_SIGNED(629,11),
TO_SIGNED(653,11),
TO_SIGNED(675,11),
TO_SIGNED(694,11),
TO_SIGNED(711,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(729,11),
TO_SIGNED(716,11),
TO_SIGNED(701,11),
TO_SIGNED(683,11),
TO_SIGNED(662,11),
TO_SIGNED(639,11),
TO_SIGNED(613,11),
TO_SIGNED(584,11),
TO_SIGNED(554,11),
TO_SIGNED(521,11),
TO_SIGNED(486,11),
TO_SIGNED(449,11),
TO_SIGNED(411,11),
TO_SIGNED(371,11),
TO_SIGNED(329,11),
TO_SIGNED(286,11),
TO_SIGNED(242,11),
TO_SIGNED(197,11),
TO_SIGNED(152,11),
TO_SIGNED(105,11),
TO_SIGNED(59,11),
TO_SIGNED(12,11),
TO_SIGNED(-35,11),
TO_SIGNED(-82,11),
TO_SIGNED(-129,11),
TO_SIGNED(-175,11),
TO_SIGNED(-220,11),
TO_SIGNED(-265,11),
TO_SIGNED(-308,11),
TO_SIGNED(-350,11),
TO_SIGNED(-391,11),
TO_SIGNED(-430,11),
TO_SIGNED(-468,11),
TO_SIGNED(-504,11),
TO_SIGNED(-538,11),
TO_SIGNED(-569,11),
TO_SIGNED(-599,11),
TO_SIGNED(-626,11),
TO_SIGNED(-651,11),
TO_SIGNED(-673,11),
TO_SIGNED(-692,11),
TO_SIGNED(-709,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-685,11),
TO_SIGNED(-664,11),
TO_SIGNED(-641,11),
TO_SIGNED(-616,11),
TO_SIGNED(-588,11),
TO_SIGNED(-557,11),
TO_SIGNED(-525,11),
TO_SIGNED(-490,11),
TO_SIGNED(-454,11),
TO_SIGNED(-415,11),
TO_SIGNED(-375,11),
TO_SIGNED(-334,11),
TO_SIGNED(-291,11),
TO_SIGNED(-247,11),
TO_SIGNED(-203,11),
TO_SIGNED(-157,11),
TO_SIGNED(-111,11),
TO_SIGNED(-64,11),
TO_SIGNED(-17,11),
TO_SIGNED(30,11),
TO_SIGNED(77,11),
TO_SIGNED(123,11),
TO_SIGNED(169,11),
TO_SIGNED(215,11),
TO_SIGNED(260,11),
TO_SIGNED(303,11),
TO_SIGNED(345,11),
TO_SIGNED(387,11),
TO_SIGNED(426,11),
TO_SIGNED(464,11),
TO_SIGNED(500,11),
TO_SIGNED(534,11),
TO_SIGNED(566,11),
TO_SIGNED(596,11),
TO_SIGNED(623,11),
TO_SIGNED(648,11),
TO_SIGNED(670,11),
TO_SIGNED(690,11),
TO_SIGNED(707,11),
TO_SIGNED(721,11),
TO_SIGNED(733,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(705,11),
TO_SIGNED(687,11),
TO_SIGNED(667,11),
TO_SIGNED(644,11),
TO_SIGNED(619,11),
TO_SIGNED(591,11),
TO_SIGNED(561,11),
TO_SIGNED(529,11),
TO_SIGNED(494,11),
TO_SIGNED(458,11),
TO_SIGNED(420,11),
TO_SIGNED(380,11),
TO_SIGNED(339,11),
TO_SIGNED(296,11),
TO_SIGNED(252,11),
TO_SIGNED(208,11),
TO_SIGNED(162,11),
TO_SIGNED(116,11),
TO_SIGNED(69,11),
TO_SIGNED(22,11),
TO_SIGNED(-25,11),
TO_SIGNED(-71,11),
TO_SIGNED(-118,11),
TO_SIGNED(-164,11),
TO_SIGNED(-210,11),
TO_SIGNED(-255,11),
TO_SIGNED(-298,11),
TO_SIGNED(-341,11),
TO_SIGNED(-382,11),
TO_SIGNED(-422,11),
TO_SIGNED(-460,11),
TO_SIGNED(-496,11),
TO_SIGNED(-530,11),
TO_SIGNED(-562,11),
TO_SIGNED(-592,11),
TO_SIGNED(-620,11),
TO_SIGNED(-645,11),
TO_SIGNED(-668,11),
TO_SIGNED(-688,11),
TO_SIGNED(-705,11),
TO_SIGNED(-720,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-721,11),
TO_SIGNED(-706,11),
TO_SIGNED(-689,11),
TO_SIGNED(-669,11),
TO_SIGNED(-647,11),
TO_SIGNED(-622,11),
TO_SIGNED(-594,11),
TO_SIGNED(-564,11),
TO_SIGNED(-532,11),
TO_SIGNED(-498,11),
TO_SIGNED(-462,11),
TO_SIGNED(-424,11),
TO_SIGNED(-385,11),
TO_SIGNED(-344,11),
TO_SIGNED(-301,11),
TO_SIGNED(-258,11),
TO_SIGNED(-213,11),
TO_SIGNED(-167,11),
TO_SIGNED(-121,11),
TO_SIGNED(-75,11),
TO_SIGNED(-28,11),
TO_SIGNED(19,11),
TO_SIGNED(66,11),
TO_SIGNED(113,11),
TO_SIGNED(159,11),
TO_SIGNED(205,11),
TO_SIGNED(249,11),
TO_SIGNED(293,11),
TO_SIGNED(336,11),
TO_SIGNED(377,11),
TO_SIGNED(417,11),
TO_SIGNED(455,11),
TO_SIGNED(492,11),
TO_SIGNED(526,11),
TO_SIGNED(559,11),
TO_SIGNED(589,11),
TO_SIGNED(617,11),
TO_SIGNED(642,11),
TO_SIGNED(665,11),
TO_SIGNED(686,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(708,11),
TO_SIGNED(691,11),
TO_SIGNED(672,11),
TO_SIGNED(650,11),
TO_SIGNED(625,11),
TO_SIGNED(598,11),
TO_SIGNED(568,11),
TO_SIGNED(536,11),
TO_SIGNED(502,11),
TO_SIGNED(466,11),
TO_SIGNED(429,11),
TO_SIGNED(389,11),
TO_SIGNED(348,11),
TO_SIGNED(306,11),
TO_SIGNED(263,11),
TO_SIGNED(218,11),
TO_SIGNED(173,11),
TO_SIGNED(127,11),
TO_SIGNED(80,11),
TO_SIGNED(33,11),
TO_SIGNED(-14,11),
TO_SIGNED(-61,11),
TO_SIGNED(-108,11),
TO_SIGNED(-154,11),
TO_SIGNED(-200,11),
TO_SIGNED(-244,11),
TO_SIGNED(-288,11),
TO_SIGNED(-331,11),
TO_SIGNED(-373,11),
TO_SIGNED(-413,11),
TO_SIGNED(-451,11),
TO_SIGNED(-488,11),
TO_SIGNED(-523,11),
TO_SIGNED(-555,11),
TO_SIGNED(-586,11),
TO_SIGNED(-614,11),
TO_SIGNED(-640,11),
TO_SIGNED(-663,11),
TO_SIGNED(-684,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-729,11),
TO_SIGNED(-739,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-710,11),
TO_SIGNED(-693,11),
TO_SIGNED(-674,11),
TO_SIGNED(-652,11),
TO_SIGNED(-628,11),
TO_SIGNED(-601,11),
TO_SIGNED(-571,11),
TO_SIGNED(-540,11),
TO_SIGNED(-506,11),
TO_SIGNED(-471,11),
TO_SIGNED(-433,11),
TO_SIGNED(-394,11),
TO_SIGNED(-353,11),
TO_SIGNED(-311,11),
TO_SIGNED(-268,11),
TO_SIGNED(-223,11),
TO_SIGNED(-178,11),
TO_SIGNED(-132,11),
TO_SIGNED(-85,11),
TO_SIGNED(-38,11),
TO_SIGNED(9,11),
TO_SIGNED(56,11),
TO_SIGNED(102,11),
TO_SIGNED(149,11),
TO_SIGNED(194,11),
TO_SIGNED(239,11),
TO_SIGNED(283,11),
TO_SIGNED(326,11),
TO_SIGNED(368,11),
TO_SIGNED(408,11),
TO_SIGNED(447,11),
TO_SIGNED(484,11),
TO_SIGNED(519,11),
TO_SIGNED(552,11),
TO_SIGNED(582,11),
TO_SIGNED(611,11),
TO_SIGNED(637,11),
TO_SIGNED(660,11),
TO_SIGNED(681,11),
TO_SIGNED(700,11),
TO_SIGNED(715,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(736,11),
TO_SIGNED(725,11),
TO_SIGNED(712,11),
TO_SIGNED(695,11),
TO_SIGNED(676,11),
TO_SIGNED(655,11),
TO_SIGNED(631,11),
TO_SIGNED(604,11),
TO_SIGNED(575,11),
TO_SIGNED(544,11),
TO_SIGNED(510,11),
TO_SIGNED(475,11),
TO_SIGNED(437,11),
TO_SIGNED(398,11),
TO_SIGNED(358,11),
TO_SIGNED(316,11),
TO_SIGNED(273,11),
TO_SIGNED(228,11),
TO_SIGNED(183,11),
TO_SIGNED(137,11),
TO_SIGNED(91,11),
TO_SIGNED(44,11),
TO_SIGNED(-3,11),
TO_SIGNED(-50,11),
TO_SIGNED(-97,11),
TO_SIGNED(-143,11),
TO_SIGNED(-189,11),
TO_SIGNED(-234,11),
TO_SIGNED(-278,11),
TO_SIGNED(-322,11),
TO_SIGNED(-363,11),
TO_SIGNED(-404,11),
TO_SIGNED(-443,11),
TO_SIGNED(-480,11),
TO_SIGNED(-515,11),
TO_SIGNED(-548,11),
TO_SIGNED(-579,11),
TO_SIGNED(-608,11),
TO_SIGNED(-634,11),
TO_SIGNED(-658,11),
TO_SIGNED(-679,11),
TO_SIGNED(-698,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-679,11),
TO_SIGNED(-657,11),
TO_SIGNED(-633,11),
TO_SIGNED(-607,11),
TO_SIGNED(-578,11),
TO_SIGNED(-547,11),
TO_SIGNED(-514,11),
TO_SIGNED(-479,11),
TO_SIGNED(-442,11),
TO_SIGNED(-403,11),
TO_SIGNED(-362,11),
TO_SIGNED(-321,11),
TO_SIGNED(-277,11),
TO_SIGNED(-233,11),
TO_SIGNED(-188,11),
TO_SIGNED(-142,11),
TO_SIGNED(-96,11),
TO_SIGNED(-49,11),
TO_SIGNED(-2,11),
TO_SIGNED(45,11),
TO_SIGNED(92,11),
TO_SIGNED(138,11),
TO_SIGNED(184,11),
TO_SIGNED(229,11),
TO_SIGNED(274,11),
TO_SIGNED(317,11),
TO_SIGNED(359,11),
TO_SIGNED(399,11),
TO_SIGNED(438,11),
TO_SIGNED(476,11),
TO_SIGNED(511,11),
TO_SIGNED(544,11),
TO_SIGNED(576,11),
TO_SIGNED(605,11),
TO_SIGNED(631,11),
TO_SIGNED(655,11),
TO_SIGNED(677,11),
TO_SIGNED(696,11),
TO_SIGNED(712,11),
TO_SIGNED(725,11),
TO_SIGNED(736,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(715,11),
TO_SIGNED(699,11),
TO_SIGNED(681,11),
TO_SIGNED(660,11),
TO_SIGNED(636,11),
TO_SIGNED(610,11),
TO_SIGNED(582,11),
TO_SIGNED(551,11),
TO_SIGNED(518,11),
TO_SIGNED(483,11),
TO_SIGNED(446,11),
TO_SIGNED(407,11),
TO_SIGNED(367,11),
TO_SIGNED(325,11),
TO_SIGNED(282,11),
TO_SIGNED(238,11),
TO_SIGNED(193,11),
TO_SIGNED(148,11),
TO_SIGNED(101,11),
TO_SIGNED(54,11),
TO_SIGNED(7,11),
TO_SIGNED(-40,11),
TO_SIGNED(-86,11),
TO_SIGNED(-133,11),
TO_SIGNED(-179,11),
TO_SIGNED(-224,11),
TO_SIGNED(-269,11),
TO_SIGNED(-312,11),
TO_SIGNED(-354,11),
TO_SIGNED(-395,11),
TO_SIGNED(-434,11),
TO_SIGNED(-471,11),
TO_SIGNED(-507,11),
TO_SIGNED(-541,11),
TO_SIGNED(-572,11),
TO_SIGNED(-601,11),
TO_SIGNED(-628,11),
TO_SIGNED(-653,11),
TO_SIGNED(-675,11),
TO_SIGNED(-694,11),
TO_SIGNED(-710,11),
TO_SIGNED(-724,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-701,11),
TO_SIGNED(-683,11),
TO_SIGNED(-662,11),
TO_SIGNED(-639,11),
TO_SIGNED(-613,11),
TO_SIGNED(-585,11),
TO_SIGNED(-554,11),
TO_SIGNED(-522,11),
TO_SIGNED(-487,11),
TO_SIGNED(-450,11),
TO_SIGNED(-412,11),
TO_SIGNED(-372,11),
TO_SIGNED(-330,11),
TO_SIGNED(-287,11),
TO_SIGNED(-243,11),
TO_SIGNED(-198,11),
TO_SIGNED(-153,11),
TO_SIGNED(-106,11),
TO_SIGNED(-60,11),
TO_SIGNED(-13,11),
TO_SIGNED(34,11),
TO_SIGNED(81,11),
TO_SIGNED(128,11),
TO_SIGNED(174,11),
TO_SIGNED(219,11),
TO_SIGNED(264,11),
TO_SIGNED(307,11),
TO_SIGNED(349,11),
TO_SIGNED(390,11),
TO_SIGNED(430,11),
TO_SIGNED(467,11),
TO_SIGNED(503,11),
TO_SIGNED(537,11),
TO_SIGNED(569,11),
TO_SIGNED(598,11),
TO_SIGNED(625,11),
TO_SIGNED(650,11),
TO_SIGNED(672,11),
TO_SIGNED(692,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(730,11),
TO_SIGNED(718,11),
TO_SIGNED(703,11),
TO_SIGNED(685,11),
TO_SIGNED(665,11),
TO_SIGNED(642,11),
TO_SIGNED(616,11),
TO_SIGNED(588,11),
TO_SIGNED(558,11),
TO_SIGNED(526,11),
TO_SIGNED(491,11),
TO_SIGNED(455,11),
TO_SIGNED(416,11),
TO_SIGNED(376,11),
TO_SIGNED(335,11),
TO_SIGNED(292,11),
TO_SIGNED(248,11),
TO_SIGNED(204,11),
TO_SIGNED(158,11),
TO_SIGNED(112,11),
TO_SIGNED(65,11),
TO_SIGNED(18,11),
TO_SIGNED(-29,11),
TO_SIGNED(-76,11),
TO_SIGNED(-122,11),
TO_SIGNED(-168,11),
TO_SIGNED(-214,11),
TO_SIGNED(-259,11),
TO_SIGNED(-302,11),
TO_SIGNED(-345,11),
TO_SIGNED(-386,11),
TO_SIGNED(-425,11),
TO_SIGNED(-463,11),
TO_SIGNED(-499,11),
TO_SIGNED(-533,11),
TO_SIGNED(-565,11),
TO_SIGNED(-595,11),
TO_SIGNED(-622,11),
TO_SIGNED(-647,11),
TO_SIGNED(-670,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-721,11),
TO_SIGNED(-733,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-720,11),
TO_SIGNED(-705,11),
TO_SIGNED(-688,11),
TO_SIGNED(-667,11),
TO_SIGNED(-645,11),
TO_SIGNED(-619,11),
TO_SIGNED(-592,11),
TO_SIGNED(-562,11),
TO_SIGNED(-529,11),
TO_SIGNED(-495,11),
TO_SIGNED(-459,11),
TO_SIGNED(-421,11),
TO_SIGNED(-381,11),
TO_SIGNED(-340,11),
TO_SIGNED(-297,11),
TO_SIGNED(-254,11),
TO_SIGNED(-209,11),
TO_SIGNED(-163,11),
TO_SIGNED(-117,11),
TO_SIGNED(-70,11),
TO_SIGNED(-24,11),
TO_SIGNED(24,11),
TO_SIGNED(70,11),
TO_SIGNED(117,11),
TO_SIGNED(163,11),
TO_SIGNED(209,11),
TO_SIGNED(254,11),
TO_SIGNED(297,11),
TO_SIGNED(340,11),
TO_SIGNED(381,11),
TO_SIGNED(421,11),
TO_SIGNED(459,11),
TO_SIGNED(495,11),
TO_SIGNED(529,11),
TO_SIGNED(562,11),
TO_SIGNED(592,11),
TO_SIGNED(619,11),
TO_SIGNED(645,11),
TO_SIGNED(667,11),
TO_SIGNED(688,11),
TO_SIGNED(705,11),
TO_SIGNED(720,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(733,11),
TO_SIGNED(721,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(670,11),
TO_SIGNED(647,11),
TO_SIGNED(622,11),
TO_SIGNED(595,11),
TO_SIGNED(565,11),
TO_SIGNED(533,11),
TO_SIGNED(499,11),
TO_SIGNED(463,11),
TO_SIGNED(425,11),
TO_SIGNED(386,11),
TO_SIGNED(345,11),
TO_SIGNED(302,11),
TO_SIGNED(259,11),
TO_SIGNED(214,11),
TO_SIGNED(168,11),
TO_SIGNED(122,11),
TO_SIGNED(76,11),
TO_SIGNED(29,11),
TO_SIGNED(-18,11),
TO_SIGNED(-65,11),
TO_SIGNED(-112,11),
TO_SIGNED(-158,11),
TO_SIGNED(-204,11),
TO_SIGNED(-248,11),
TO_SIGNED(-292,11),
TO_SIGNED(-335,11),
TO_SIGNED(-376,11),
TO_SIGNED(-416,11),
TO_SIGNED(-455,11),
TO_SIGNED(-491,11),
TO_SIGNED(-526,11),
TO_SIGNED(-558,11),
TO_SIGNED(-588,11),
TO_SIGNED(-616,11),
TO_SIGNED(-642,11),
TO_SIGNED(-665,11),
TO_SIGNED(-685,11),
TO_SIGNED(-703,11),
TO_SIGNED(-718,11),
TO_SIGNED(-730,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-692,11),
TO_SIGNED(-672,11),
TO_SIGNED(-650,11),
TO_SIGNED(-625,11),
TO_SIGNED(-598,11),
TO_SIGNED(-569,11),
TO_SIGNED(-537,11),
TO_SIGNED(-503,11),
TO_SIGNED(-467,11),
TO_SIGNED(-430,11),
TO_SIGNED(-390,11),
TO_SIGNED(-349,11),
TO_SIGNED(-307,11),
TO_SIGNED(-264,11),
TO_SIGNED(-219,11),
TO_SIGNED(-174,11),
TO_SIGNED(-128,11),
TO_SIGNED(-81,11),
TO_SIGNED(-34,11),
TO_SIGNED(13,11),
TO_SIGNED(60,11),
TO_SIGNED(106,11),
TO_SIGNED(153,11),
TO_SIGNED(198,11),
TO_SIGNED(243,11),
TO_SIGNED(287,11),
TO_SIGNED(330,11),
TO_SIGNED(372,11),
TO_SIGNED(412,11),
TO_SIGNED(450,11),
TO_SIGNED(487,11),
TO_SIGNED(522,11),
TO_SIGNED(554,11),
TO_SIGNED(585,11),
TO_SIGNED(613,11),
TO_SIGNED(639,11),
TO_SIGNED(662,11),
TO_SIGNED(683,11),
TO_SIGNED(701,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(724,11),
TO_SIGNED(710,11),
TO_SIGNED(694,11),
TO_SIGNED(675,11),
TO_SIGNED(653,11),
TO_SIGNED(628,11),
TO_SIGNED(601,11),
TO_SIGNED(572,11),
TO_SIGNED(541,11),
TO_SIGNED(507,11),
TO_SIGNED(471,11),
TO_SIGNED(434,11),
TO_SIGNED(395,11),
TO_SIGNED(354,11),
TO_SIGNED(312,11),
TO_SIGNED(269,11),
TO_SIGNED(224,11),
TO_SIGNED(179,11),
TO_SIGNED(133,11),
TO_SIGNED(86,11),
TO_SIGNED(40,11),
TO_SIGNED(-7,11),
TO_SIGNED(-54,11),
TO_SIGNED(-101,11),
TO_SIGNED(-148,11),
TO_SIGNED(-193,11),
TO_SIGNED(-238,11),
TO_SIGNED(-282,11),
TO_SIGNED(-325,11),
TO_SIGNED(-367,11),
TO_SIGNED(-407,11),
TO_SIGNED(-446,11),
TO_SIGNED(-483,11),
TO_SIGNED(-518,11),
TO_SIGNED(-551,11),
TO_SIGNED(-582,11),
TO_SIGNED(-610,11),
TO_SIGNED(-636,11),
TO_SIGNED(-660,11),
TO_SIGNED(-681,11),
TO_SIGNED(-699,11),
TO_SIGNED(-715,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-736,11),
TO_SIGNED(-725,11),
TO_SIGNED(-712,11),
TO_SIGNED(-696,11),
TO_SIGNED(-677,11),
TO_SIGNED(-655,11),
TO_SIGNED(-631,11),
TO_SIGNED(-605,11),
TO_SIGNED(-576,11),
TO_SIGNED(-544,11),
TO_SIGNED(-511,11),
TO_SIGNED(-476,11),
TO_SIGNED(-438,11),
TO_SIGNED(-399,11),
TO_SIGNED(-359,11),
TO_SIGNED(-317,11),
TO_SIGNED(-274,11),
TO_SIGNED(-229,11),
TO_SIGNED(-184,11),
TO_SIGNED(-138,11),
TO_SIGNED(-92,11),
TO_SIGNED(-45,11),
TO_SIGNED(2,11),
TO_SIGNED(49,11),
TO_SIGNED(96,11),
TO_SIGNED(142,11),
TO_SIGNED(188,11),
TO_SIGNED(233,11),
TO_SIGNED(277,11),
TO_SIGNED(321,11),
TO_SIGNED(362,11),
TO_SIGNED(403,11),
TO_SIGNED(442,11),
TO_SIGNED(479,11),
TO_SIGNED(514,11),
TO_SIGNED(547,11),
TO_SIGNED(578,11),
TO_SIGNED(607,11),
TO_SIGNED(633,11),
TO_SIGNED(657,11),
TO_SIGNED(679,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(698,11),
TO_SIGNED(679,11),
TO_SIGNED(658,11),
TO_SIGNED(634,11),
TO_SIGNED(608,11),
TO_SIGNED(579,11),
TO_SIGNED(548,11),
TO_SIGNED(515,11),
TO_SIGNED(480,11),
TO_SIGNED(443,11),
TO_SIGNED(404,11),
TO_SIGNED(363,11),
TO_SIGNED(322,11),
TO_SIGNED(278,11),
TO_SIGNED(234,11),
TO_SIGNED(189,11),
TO_SIGNED(143,11),
TO_SIGNED(97,11),
TO_SIGNED(50,11),
TO_SIGNED(3,11),
TO_SIGNED(-44,11),
TO_SIGNED(-91,11),
TO_SIGNED(-137,11),
TO_SIGNED(-183,11),
TO_SIGNED(-228,11),
TO_SIGNED(-273,11),
TO_SIGNED(-316,11),
TO_SIGNED(-358,11),
TO_SIGNED(-398,11),
TO_SIGNED(-437,11),
TO_SIGNED(-475,11),
TO_SIGNED(-510,11),
TO_SIGNED(-544,11),
TO_SIGNED(-575,11),
TO_SIGNED(-604,11),
TO_SIGNED(-631,11),
TO_SIGNED(-655,11),
TO_SIGNED(-676,11),
TO_SIGNED(-695,11),
TO_SIGNED(-712,11),
TO_SIGNED(-725,11),
TO_SIGNED(-736,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-715,11),
TO_SIGNED(-700,11),
TO_SIGNED(-681,11),
TO_SIGNED(-660,11),
TO_SIGNED(-637,11),
TO_SIGNED(-611,11),
TO_SIGNED(-582,11),
TO_SIGNED(-552,11),
TO_SIGNED(-519,11),
TO_SIGNED(-484,11),
TO_SIGNED(-447,11),
TO_SIGNED(-408,11),
TO_SIGNED(-368,11),
TO_SIGNED(-326,11),
TO_SIGNED(-283,11),
TO_SIGNED(-239,11),
TO_SIGNED(-194,11),
TO_SIGNED(-149,11),
TO_SIGNED(-102,11),
TO_SIGNED(-56,11),
TO_SIGNED(-9,11),
TO_SIGNED(38,11),
TO_SIGNED(85,11),
TO_SIGNED(132,11),
TO_SIGNED(178,11),
TO_SIGNED(223,11),
TO_SIGNED(268,11),
TO_SIGNED(311,11),
TO_SIGNED(353,11),
TO_SIGNED(394,11),
TO_SIGNED(433,11),
TO_SIGNED(471,11),
TO_SIGNED(506,11),
TO_SIGNED(540,11),
TO_SIGNED(571,11),
TO_SIGNED(601,11),
TO_SIGNED(628,11),
TO_SIGNED(652,11),
TO_SIGNED(674,11),
TO_SIGNED(693,11),
TO_SIGNED(710,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(739,11),
TO_SIGNED(729,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(684,11),
TO_SIGNED(663,11),
TO_SIGNED(640,11),
TO_SIGNED(614,11),
TO_SIGNED(586,11),
TO_SIGNED(555,11),
TO_SIGNED(523,11),
TO_SIGNED(488,11),
TO_SIGNED(451,11),
TO_SIGNED(413,11),
TO_SIGNED(373,11),
TO_SIGNED(331,11),
TO_SIGNED(288,11),
TO_SIGNED(244,11),
TO_SIGNED(200,11),
TO_SIGNED(154,11),
TO_SIGNED(108,11),
TO_SIGNED(61,11),
TO_SIGNED(14,11),
TO_SIGNED(-33,11),
TO_SIGNED(-80,11),
TO_SIGNED(-127,11),
TO_SIGNED(-173,11),
TO_SIGNED(-218,11),
TO_SIGNED(-263,11),
TO_SIGNED(-306,11),
TO_SIGNED(-348,11),
TO_SIGNED(-389,11),
TO_SIGNED(-429,11),
TO_SIGNED(-466,11),
TO_SIGNED(-502,11),
TO_SIGNED(-536,11),
TO_SIGNED(-568,11),
TO_SIGNED(-598,11),
TO_SIGNED(-625,11),
TO_SIGNED(-650,11),
TO_SIGNED(-672,11),
TO_SIGNED(-691,11),
TO_SIGNED(-708,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-686,11),
TO_SIGNED(-665,11),
TO_SIGNED(-642,11),
TO_SIGNED(-617,11),
TO_SIGNED(-589,11),
TO_SIGNED(-559,11),
TO_SIGNED(-526,11),
TO_SIGNED(-492,11),
TO_SIGNED(-455,11),
TO_SIGNED(-417,11),
TO_SIGNED(-377,11),
TO_SIGNED(-336,11),
TO_SIGNED(-293,11),
TO_SIGNED(-249,11),
TO_SIGNED(-205,11),
TO_SIGNED(-159,11),
TO_SIGNED(-113,11),
TO_SIGNED(-66,11),
TO_SIGNED(-19,11),
TO_SIGNED(28,11),
TO_SIGNED(75,11),
TO_SIGNED(121,11),
TO_SIGNED(167,11),
TO_SIGNED(213,11),
TO_SIGNED(258,11),
TO_SIGNED(301,11),
TO_SIGNED(344,11),
TO_SIGNED(385,11),
TO_SIGNED(424,11),
TO_SIGNED(462,11),
TO_SIGNED(498,11),
TO_SIGNED(532,11),
TO_SIGNED(564,11),
TO_SIGNED(594,11),
TO_SIGNED(622,11),
TO_SIGNED(647,11),
TO_SIGNED(669,11),
TO_SIGNED(689,11),
TO_SIGNED(706,11),
TO_SIGNED(721,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(720,11),
TO_SIGNED(705,11),
TO_SIGNED(688,11),
TO_SIGNED(668,11),
TO_SIGNED(645,11),
TO_SIGNED(620,11),
TO_SIGNED(592,11),
TO_SIGNED(562,11),
TO_SIGNED(530,11),
TO_SIGNED(496,11),
TO_SIGNED(460,11),
TO_SIGNED(422,11),
TO_SIGNED(382,11),
TO_SIGNED(341,11),
TO_SIGNED(298,11),
TO_SIGNED(255,11),
TO_SIGNED(210,11),
TO_SIGNED(164,11),
TO_SIGNED(118,11),
TO_SIGNED(71,11),
TO_SIGNED(25,11),
TO_SIGNED(-22,11),
TO_SIGNED(-69,11),
TO_SIGNED(-116,11),
TO_SIGNED(-162,11),
TO_SIGNED(-208,11),
TO_SIGNED(-252,11),
TO_SIGNED(-296,11),
TO_SIGNED(-339,11),
TO_SIGNED(-380,11),
TO_SIGNED(-420,11),
TO_SIGNED(-458,11),
TO_SIGNED(-494,11),
TO_SIGNED(-529,11),
TO_SIGNED(-561,11),
TO_SIGNED(-591,11),
TO_SIGNED(-619,11),
TO_SIGNED(-644,11),
TO_SIGNED(-667,11),
TO_SIGNED(-687,11),
TO_SIGNED(-705,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-733,11),
TO_SIGNED(-721,11),
TO_SIGNED(-707,11),
TO_SIGNED(-690,11),
TO_SIGNED(-670,11),
TO_SIGNED(-648,11),
TO_SIGNED(-623,11),
TO_SIGNED(-596,11),
TO_SIGNED(-566,11),
TO_SIGNED(-534,11),
TO_SIGNED(-500,11),
TO_SIGNED(-464,11),
TO_SIGNED(-426,11),
TO_SIGNED(-387,11),
TO_SIGNED(-345,11),
TO_SIGNED(-303,11),
TO_SIGNED(-260,11),
TO_SIGNED(-215,11),
TO_SIGNED(-169,11),
TO_SIGNED(-123,11),
TO_SIGNED(-77,11),
TO_SIGNED(-30,11),
TO_SIGNED(17,11),
TO_SIGNED(64,11),
TO_SIGNED(111,11),
TO_SIGNED(157,11),
TO_SIGNED(203,11),
TO_SIGNED(247,11),
TO_SIGNED(291,11),
TO_SIGNED(334,11),
TO_SIGNED(375,11),
TO_SIGNED(415,11),
TO_SIGNED(454,11),
TO_SIGNED(490,11),
TO_SIGNED(525,11),
TO_SIGNED(557,11),
TO_SIGNED(588,11),
TO_SIGNED(616,11),
TO_SIGNED(641,11),
TO_SIGNED(664,11),
TO_SIGNED(685,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(709,11),
TO_SIGNED(692,11),
TO_SIGNED(673,11),
TO_SIGNED(651,11),
TO_SIGNED(626,11),
TO_SIGNED(599,11),
TO_SIGNED(569,11),
TO_SIGNED(538,11),
TO_SIGNED(504,11),
TO_SIGNED(468,11),
TO_SIGNED(430,11),
TO_SIGNED(391,11),
TO_SIGNED(350,11),
TO_SIGNED(308,11),
TO_SIGNED(265,11),
TO_SIGNED(220,11),
TO_SIGNED(175,11),
TO_SIGNED(129,11),
TO_SIGNED(82,11),
TO_SIGNED(35,11),
TO_SIGNED(-12,11),
TO_SIGNED(-59,11),
TO_SIGNED(-105,11),
TO_SIGNED(-152,11),
TO_SIGNED(-197,11),
TO_SIGNED(-242,11),
TO_SIGNED(-286,11),
TO_SIGNED(-329,11),
TO_SIGNED(-371,11),
TO_SIGNED(-411,11),
TO_SIGNED(-449,11),
TO_SIGNED(-486,11),
TO_SIGNED(-521,11),
TO_SIGNED(-554,11),
TO_SIGNED(-584,11),
TO_SIGNED(-613,11),
TO_SIGNED(-639,11),
TO_SIGNED(-662,11),
TO_SIGNED(-683,11),
TO_SIGNED(-701,11),
TO_SIGNED(-716,11),
TO_SIGNED(-729,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-711,11),
TO_SIGNED(-694,11),
TO_SIGNED(-675,11),
TO_SIGNED(-653,11),
TO_SIGNED(-629,11),
TO_SIGNED(-602,11),
TO_SIGNED(-573,11),
TO_SIGNED(-541,11),
TO_SIGNED(-508,11),
TO_SIGNED(-472,11),
TO_SIGNED(-435,11),
TO_SIGNED(-396,11),
TO_SIGNED(-355,11),
TO_SIGNED(-313,11),
TO_SIGNED(-270,11),
TO_SIGNED(-225,11),
TO_SIGNED(-180,11),
TO_SIGNED(-134,11),
TO_SIGNED(-87,11),
TO_SIGNED(-41,11),
TO_SIGNED(6,11),
TO_SIGNED(53,11),
TO_SIGNED(100,11),
TO_SIGNED(147,11),
TO_SIGNED(192,11),
TO_SIGNED(237,11),
TO_SIGNED(281,11),
TO_SIGNED(324,11),
TO_SIGNED(366,11),
TO_SIGNED(406,11),
TO_SIGNED(445,11),
TO_SIGNED(482,11),
TO_SIGNED(517,11),
TO_SIGNED(550,11),
TO_SIGNED(581,11),
TO_SIGNED(610,11),
TO_SIGNED(636,11),
TO_SIGNED(659,11),
TO_SIGNED(681,11),
TO_SIGNED(699,11),
TO_SIGNED(715,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(712,11),
TO_SIGNED(696,11),
TO_SIGNED(677,11),
TO_SIGNED(656,11),
TO_SIGNED(632,11),
TO_SIGNED(605,11),
TO_SIGNED(576,11),
TO_SIGNED(545,11),
TO_SIGNED(512,11),
TO_SIGNED(476,11),
TO_SIGNED(439,11),
TO_SIGNED(400,11),
TO_SIGNED(360,11),
TO_SIGNED(318,11),
TO_SIGNED(275,11),
TO_SIGNED(230,11),
TO_SIGNED(185,11),
TO_SIGNED(139,11),
TO_SIGNED(93,11),
TO_SIGNED(46,11),
TO_SIGNED(-1,11),
TO_SIGNED(-48,11),
TO_SIGNED(-95,11),
TO_SIGNED(-141,11),
TO_SIGNED(-187,11),
TO_SIGNED(-232,11),
TO_SIGNED(-276,11),
TO_SIGNED(-320,11),
TO_SIGNED(-362,11),
TO_SIGNED(-402,11),
TO_SIGNED(-441,11),
TO_SIGNED(-478,11),
TO_SIGNED(-513,11),
TO_SIGNED(-547,11),
TO_SIGNED(-578,11),
TO_SIGNED(-606,11),
TO_SIGNED(-633,11),
TO_SIGNED(-657,11),
TO_SIGNED(-678,11),
TO_SIGNED(-697,11),
TO_SIGNED(-713,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-714,11),
TO_SIGNED(-698,11),
TO_SIGNED(-680,11),
TO_SIGNED(-658,11),
TO_SIGNED(-635,11),
TO_SIGNED(-608,11),
TO_SIGNED(-580,11),
TO_SIGNED(-549,11),
TO_SIGNED(-516,11),
TO_SIGNED(-480,11),
TO_SIGNED(-443,11),
TO_SIGNED(-405,11),
TO_SIGNED(-364,11),
TO_SIGNED(-323,11),
TO_SIGNED(-279,11),
TO_SIGNED(-235,11),
TO_SIGNED(-190,11),
TO_SIGNED(-144,11),
TO_SIGNED(-98,11),
TO_SIGNED(-51,11),
TO_SIGNED(-4,11),
TO_SIGNED(43,11),
TO_SIGNED(90,11),
TO_SIGNED(136,11),
TO_SIGNED(182,11),
TO_SIGNED(227,11),
TO_SIGNED(272,11),
TO_SIGNED(315,11),
TO_SIGNED(357,11),
TO_SIGNED(397,11),
TO_SIGNED(437,11),
TO_SIGNED(474,11),
TO_SIGNED(509,11),
TO_SIGNED(543,11),
TO_SIGNED(574,11),
TO_SIGNED(603,11),
TO_SIGNED(630,11),
TO_SIGNED(654,11),
TO_SIGNED(676,11),
TO_SIGNED(695,11),
TO_SIGNED(711,11),
TO_SIGNED(725,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(716,11),
TO_SIGNED(700,11),
TO_SIGNED(682,11),
TO_SIGNED(661,11),
TO_SIGNED(637,11),
TO_SIGNED(611,11),
TO_SIGNED(583,11),
TO_SIGNED(552,11),
TO_SIGNED(519,11),
TO_SIGNED(485,11),
TO_SIGNED(448,11),
TO_SIGNED(409,11),
TO_SIGNED(369,11),
TO_SIGNED(327,11),
TO_SIGNED(284,11),
TO_SIGNED(240,11),
TO_SIGNED(195,11),
TO_SIGNED(150,11),
TO_SIGNED(103,11),
TO_SIGNED(57,11),
TO_SIGNED(10,11),
TO_SIGNED(-37,11),
TO_SIGNED(-84,11),
TO_SIGNED(-131,11),
TO_SIGNED(-177,11),
TO_SIGNED(-222,11),
TO_SIGNED(-267,11),
TO_SIGNED(-310,11),
TO_SIGNED(-352,11),
TO_SIGNED(-393,11),
TO_SIGNED(-432,11),
TO_SIGNED(-470,11),
TO_SIGNED(-505,11),
TO_SIGNED(-539,11),
TO_SIGNED(-571,11),
TO_SIGNED(-600,11),
TO_SIGNED(-627,11),
TO_SIGNED(-652,11),
TO_SIGNED(-674,11),
TO_SIGNED(-693,11),
TO_SIGNED(-710,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-702,11),
TO_SIGNED(-684,11),
TO_SIGNED(-663,11),
TO_SIGNED(-640,11),
TO_SIGNED(-615,11),
TO_SIGNED(-586,11),
TO_SIGNED(-556,11),
TO_SIGNED(-523,11),
TO_SIGNED(-489,11),
TO_SIGNED(-452,11),
TO_SIGNED(-414,11),
TO_SIGNED(-374,11),
TO_SIGNED(-332,11),
TO_SIGNED(-289,11),
TO_SIGNED(-245,11),
TO_SIGNED(-201,11),
TO_SIGNED(-155,11),
TO_SIGNED(-109,11),
TO_SIGNED(-62,11),
TO_SIGNED(-15,11),
TO_SIGNED(32,11),
TO_SIGNED(79,11),
TO_SIGNED(125,11),
TO_SIGNED(172,11),
TO_SIGNED(217,11),
TO_SIGNED(262,11),
TO_SIGNED(305,11),
TO_SIGNED(347,11),
TO_SIGNED(388,11),
TO_SIGNED(428,11),
TO_SIGNED(466,11),
TO_SIGNED(501,11),
TO_SIGNED(535,11),
TO_SIGNED(567,11),
TO_SIGNED(597,11),
TO_SIGNED(624,11),
TO_SIGNED(649,11),
TO_SIGNED(671,11),
TO_SIGNED(691,11),
TO_SIGNED(708,11),
TO_SIGNED(722,11),
TO_SIGNED(733,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(704,11),
TO_SIGNED(686,11),
TO_SIGNED(666,11),
TO_SIGNED(643,11),
TO_SIGNED(618,11),
TO_SIGNED(590,11),
TO_SIGNED(559,11),
TO_SIGNED(527,11),
TO_SIGNED(493,11),
TO_SIGNED(456,11),
TO_SIGNED(418,11),
TO_SIGNED(378,11),
TO_SIGNED(337,11),
TO_SIGNED(294,11),
TO_SIGNED(250,11),
TO_SIGNED(206,11),
TO_SIGNED(160,11),
TO_SIGNED(114,11),
TO_SIGNED(67,11),
TO_SIGNED(20,11),
TO_SIGNED(-27,11),
TO_SIGNED(-74,11),
TO_SIGNED(-120,11),
TO_SIGNED(-166,11),
TO_SIGNED(-212,11),
TO_SIGNED(-257,11),
TO_SIGNED(-300,11),
TO_SIGNED(-343,11),
TO_SIGNED(-384,11),
TO_SIGNED(-423,11),
TO_SIGNED(-461,11),
TO_SIGNED(-497,11),
TO_SIGNED(-532,11),
TO_SIGNED(-564,11),
TO_SIGNED(-594,11),
TO_SIGNED(-621,11),
TO_SIGNED(-646,11),
TO_SIGNED(-669,11),
TO_SIGNED(-689,11),
TO_SIGNED(-706,11),
TO_SIGNED(-721,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-720,11),
TO_SIGNED(-706,11),
TO_SIGNED(-688,11),
TO_SIGNED(-668,11),
TO_SIGNED(-646,11),
TO_SIGNED(-621,11),
TO_SIGNED(-593,11),
TO_SIGNED(-563,11),
TO_SIGNED(-531,11),
TO_SIGNED(-497,11),
TO_SIGNED(-460,11),
TO_SIGNED(-422,11),
TO_SIGNED(-383,11),
TO_SIGNED(-342,11),
TO_SIGNED(-299,11),
TO_SIGNED(-256,11),
TO_SIGNED(-211,11),
TO_SIGNED(-165,11),
TO_SIGNED(-119,11),
TO_SIGNED(-73,11),
TO_SIGNED(-26,11),
TO_SIGNED(21,11),
TO_SIGNED(68,11),
TO_SIGNED(115,11),
TO_SIGNED(161,11),
TO_SIGNED(207,11),
TO_SIGNED(251,11),
TO_SIGNED(295,11),
TO_SIGNED(338,11),
TO_SIGNED(379,11),
TO_SIGNED(419,11),
TO_SIGNED(457,11),
TO_SIGNED(493,11),
TO_SIGNED(528,11),
TO_SIGNED(560,11),
TO_SIGNED(590,11),
TO_SIGNED(618,11),
TO_SIGNED(644,11),
TO_SIGNED(666,11),
TO_SIGNED(687,11),
TO_SIGNED(704,11),
TO_SIGNED(719,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(671,11),
TO_SIGNED(648,11),
TO_SIGNED(624,11),
TO_SIGNED(596,11),
TO_SIGNED(567,11),
TO_SIGNED(535,11),
TO_SIGNED(501,11),
TO_SIGNED(465,11),
TO_SIGNED(427,11),
TO_SIGNED(387,11),
TO_SIGNED(346,11),
TO_SIGNED(304,11),
TO_SIGNED(261,11),
TO_SIGNED(216,11),
TO_SIGNED(171,11),
TO_SIGNED(124,11),
TO_SIGNED(78,11),
TO_SIGNED(31,11),
TO_SIGNED(-16,11),
TO_SIGNED(-63,11),
TO_SIGNED(-110,11),
TO_SIGNED(-156,11),
TO_SIGNED(-202,11),
TO_SIGNED(-246,11),
TO_SIGNED(-290,11),
TO_SIGNED(-333,11),
TO_SIGNED(-375,11),
TO_SIGNED(-415,11),
TO_SIGNED(-453,11),
TO_SIGNED(-489,11),
TO_SIGNED(-524,11),
TO_SIGNED(-557,11),
TO_SIGNED(-587,11),
TO_SIGNED(-615,11),
TO_SIGNED(-641,11),
TO_SIGNED(-664,11),
TO_SIGNED(-685,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-730,11),
TO_SIGNED(-739,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-693,11),
TO_SIGNED(-673,11),
TO_SIGNED(-651,11),
TO_SIGNED(-627,11),
TO_SIGNED(-599,11),
TO_SIGNED(-570,11),
TO_SIGNED(-538,11),
TO_SIGNED(-505,11),
TO_SIGNED(-469,11),
TO_SIGNED(-431,11),
TO_SIGNED(-392,11),
TO_SIGNED(-351,11),
TO_SIGNED(-309,11),
TO_SIGNED(-266,11),
TO_SIGNED(-221,11),
TO_SIGNED(-176,11),
TO_SIGNED(-130,11),
TO_SIGNED(-83,11),
TO_SIGNED(-36,11),
TO_SIGNED(11,11),
TO_SIGNED(58,11),
TO_SIGNED(104,11),
TO_SIGNED(151,11),
TO_SIGNED(196,11),
TO_SIGNED(241,11),
TO_SIGNED(285,11),
TO_SIGNED(328,11),
TO_SIGNED(370,11),
TO_SIGNED(410,11),
TO_SIGNED(449,11),
TO_SIGNED(485,11),
TO_SIGNED(520,11),
TO_SIGNED(553,11),
TO_SIGNED(584,11),
TO_SIGNED(612,11),
TO_SIGNED(638,11),
TO_SIGNED(661,11),
TO_SIGNED(682,11),
TO_SIGNED(700,11),
TO_SIGNED(716,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(725,11),
TO_SIGNED(711,11),
TO_SIGNED(695,11),
TO_SIGNED(675,11),
TO_SIGNED(654,11),
TO_SIGNED(629,11),
TO_SIGNED(603,11),
TO_SIGNED(574,11),
TO_SIGNED(542,11),
TO_SIGNED(509,11),
TO_SIGNED(473,11),
TO_SIGNED(436,11),
TO_SIGNED(397,11),
TO_SIGNED(356,11),
TO_SIGNED(314,11),
TO_SIGNED(271,11),
TO_SIGNED(226,11),
TO_SIGNED(181,11),
TO_SIGNED(135,11),
TO_SIGNED(88,11),
TO_SIGNED(42,11),
TO_SIGNED(-5,11),
TO_SIGNED(-52,11),
TO_SIGNED(-99,11),
TO_SIGNED(-145,11),
TO_SIGNED(-191,11),
TO_SIGNED(-236,11),
TO_SIGNED(-280,11),
TO_SIGNED(-323,11),
TO_SIGNED(-365,11),
TO_SIGNED(-406,11),
TO_SIGNED(-444,11),
TO_SIGNED(-481,11),
TO_SIGNED(-516,11),
TO_SIGNED(-549,11),
TO_SIGNED(-580,11),
TO_SIGNED(-609,11),
TO_SIGNED(-635,11),
TO_SIGNED(-659,11),
TO_SIGNED(-680,11),
TO_SIGNED(-699,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-736,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-678,11),
TO_SIGNED(-656,11),
TO_SIGNED(-632,11),
TO_SIGNED(-606,11),
TO_SIGNED(-577,11),
TO_SIGNED(-546,11),
TO_SIGNED(-512,11),
TO_SIGNED(-477,11),
TO_SIGNED(-440,11),
TO_SIGNED(-401,11),
TO_SIGNED(-361,11),
TO_SIGNED(-319,11),
TO_SIGNED(-275,11),
TO_SIGNED(-231,11),
TO_SIGNED(-186,11),
TO_SIGNED(-140,11),
TO_SIGNED(-94,11),
TO_SIGNED(-47,11),
TO_SIGNED(0,11),
TO_SIGNED(47,11),
TO_SIGNED(94,11),
TO_SIGNED(140,11),
TO_SIGNED(186,11),
TO_SIGNED(231,11),
TO_SIGNED(275,11),
TO_SIGNED(319,11),
TO_SIGNED(361,11),
TO_SIGNED(401,11),
TO_SIGNED(440,11),
TO_SIGNED(477,11),
TO_SIGNED(512,11),
TO_SIGNED(546,11),
TO_SIGNED(577,11),
TO_SIGNED(606,11),
TO_SIGNED(632,11),
TO_SIGNED(656,11),
TO_SIGNED(678,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(736,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(699,11),
TO_SIGNED(680,11),
TO_SIGNED(659,11),
TO_SIGNED(635,11),
TO_SIGNED(609,11),
TO_SIGNED(580,11),
TO_SIGNED(549,11),
TO_SIGNED(516,11),
TO_SIGNED(481,11),
TO_SIGNED(444,11),
TO_SIGNED(406,11),
TO_SIGNED(365,11),
TO_SIGNED(323,11),
TO_SIGNED(280,11),
TO_SIGNED(236,11),
TO_SIGNED(191,11),
TO_SIGNED(145,11),
TO_SIGNED(99,11),
TO_SIGNED(52,11),
TO_SIGNED(5,11),
TO_SIGNED(-42,11),
TO_SIGNED(-88,11),
TO_SIGNED(-135,11),
TO_SIGNED(-181,11),
TO_SIGNED(-226,11),
TO_SIGNED(-271,11),
TO_SIGNED(-314,11),
TO_SIGNED(-356,11),
TO_SIGNED(-397,11),
TO_SIGNED(-436,11),
TO_SIGNED(-473,11),
TO_SIGNED(-509,11),
TO_SIGNED(-542,11),
TO_SIGNED(-574,11),
TO_SIGNED(-603,11),
TO_SIGNED(-629,11),
TO_SIGNED(-654,11),
TO_SIGNED(-675,11),
TO_SIGNED(-695,11),
TO_SIGNED(-711,11),
TO_SIGNED(-725,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-716,11),
TO_SIGNED(-700,11),
TO_SIGNED(-682,11),
TO_SIGNED(-661,11),
TO_SIGNED(-638,11),
TO_SIGNED(-612,11),
TO_SIGNED(-584,11),
TO_SIGNED(-553,11),
TO_SIGNED(-520,11),
TO_SIGNED(-485,11),
TO_SIGNED(-449,11),
TO_SIGNED(-410,11),
TO_SIGNED(-370,11),
TO_SIGNED(-328,11),
TO_SIGNED(-285,11),
TO_SIGNED(-241,11),
TO_SIGNED(-196,11),
TO_SIGNED(-151,11),
TO_SIGNED(-104,11),
TO_SIGNED(-58,11),
TO_SIGNED(-11,11),
TO_SIGNED(36,11),
TO_SIGNED(83,11),
TO_SIGNED(130,11),
TO_SIGNED(176,11),
TO_SIGNED(221,11),
TO_SIGNED(266,11),
TO_SIGNED(309,11),
TO_SIGNED(351,11),
TO_SIGNED(392,11),
TO_SIGNED(431,11),
TO_SIGNED(469,11),
TO_SIGNED(505,11),
TO_SIGNED(538,11),
TO_SIGNED(570,11),
TO_SIGNED(599,11),
TO_SIGNED(627,11),
TO_SIGNED(651,11),
TO_SIGNED(673,11),
TO_SIGNED(693,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(739,11),
TO_SIGNED(730,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(685,11),
TO_SIGNED(664,11),
TO_SIGNED(641,11),
TO_SIGNED(615,11),
TO_SIGNED(587,11),
TO_SIGNED(557,11),
TO_SIGNED(524,11),
TO_SIGNED(489,11),
TO_SIGNED(453,11),
TO_SIGNED(415,11),
TO_SIGNED(375,11),
TO_SIGNED(333,11),
TO_SIGNED(290,11),
TO_SIGNED(246,11),
TO_SIGNED(202,11),
TO_SIGNED(156,11),
TO_SIGNED(110,11),
TO_SIGNED(63,11),
TO_SIGNED(16,11),
TO_SIGNED(-31,11),
TO_SIGNED(-78,11),
TO_SIGNED(-124,11),
TO_SIGNED(-171,11),
TO_SIGNED(-216,11),
TO_SIGNED(-261,11),
TO_SIGNED(-304,11),
TO_SIGNED(-346,11),
TO_SIGNED(-387,11),
TO_SIGNED(-427,11),
TO_SIGNED(-465,11),
TO_SIGNED(-501,11),
TO_SIGNED(-535,11),
TO_SIGNED(-567,11),
TO_SIGNED(-596,11),
TO_SIGNED(-624,11),
TO_SIGNED(-648,11),
TO_SIGNED(-671,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-719,11),
TO_SIGNED(-704,11),
TO_SIGNED(-687,11),
TO_SIGNED(-666,11),
TO_SIGNED(-644,11),
TO_SIGNED(-618,11),
TO_SIGNED(-590,11),
TO_SIGNED(-560,11),
TO_SIGNED(-528,11),
TO_SIGNED(-493,11),
TO_SIGNED(-457,11),
TO_SIGNED(-419,11),
TO_SIGNED(-379,11),
TO_SIGNED(-338,11),
TO_SIGNED(-295,11),
TO_SIGNED(-251,11),
TO_SIGNED(-207,11),
TO_SIGNED(-161,11),
TO_SIGNED(-115,11),
TO_SIGNED(-68,11),
TO_SIGNED(-21,11),
TO_SIGNED(26,11),
TO_SIGNED(73,11),
TO_SIGNED(119,11),
TO_SIGNED(165,11),
TO_SIGNED(211,11),
TO_SIGNED(256,11),
TO_SIGNED(299,11),
TO_SIGNED(342,11),
TO_SIGNED(383,11),
TO_SIGNED(422,11),
TO_SIGNED(460,11),
TO_SIGNED(497,11),
TO_SIGNED(531,11),
TO_SIGNED(563,11),
TO_SIGNED(593,11),
TO_SIGNED(621,11),
TO_SIGNED(646,11),
TO_SIGNED(668,11),
TO_SIGNED(688,11),
TO_SIGNED(706,11),
TO_SIGNED(720,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(721,11),
TO_SIGNED(706,11),
TO_SIGNED(689,11),
TO_SIGNED(669,11),
TO_SIGNED(646,11),
TO_SIGNED(621,11),
TO_SIGNED(594,11),
TO_SIGNED(564,11),
TO_SIGNED(532,11),
TO_SIGNED(497,11),
TO_SIGNED(461,11),
TO_SIGNED(423,11),
TO_SIGNED(384,11),
TO_SIGNED(343,11),
TO_SIGNED(300,11),
TO_SIGNED(257,11),
TO_SIGNED(212,11),
TO_SIGNED(166,11),
TO_SIGNED(120,11),
TO_SIGNED(74,11),
TO_SIGNED(27,11),
TO_SIGNED(-20,11),
TO_SIGNED(-67,11),
TO_SIGNED(-114,11),
TO_SIGNED(-160,11),
TO_SIGNED(-206,11),
TO_SIGNED(-250,11),
TO_SIGNED(-294,11),
TO_SIGNED(-337,11),
TO_SIGNED(-378,11),
TO_SIGNED(-418,11),
TO_SIGNED(-456,11),
TO_SIGNED(-493,11),
TO_SIGNED(-527,11),
TO_SIGNED(-559,11),
TO_SIGNED(-590,11),
TO_SIGNED(-618,11),
TO_SIGNED(-643,11),
TO_SIGNED(-666,11),
TO_SIGNED(-686,11),
TO_SIGNED(-704,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-733,11),
TO_SIGNED(-722,11),
TO_SIGNED(-708,11),
TO_SIGNED(-691,11),
TO_SIGNED(-671,11),
TO_SIGNED(-649,11),
TO_SIGNED(-624,11),
TO_SIGNED(-597,11),
TO_SIGNED(-567,11),
TO_SIGNED(-535,11),
TO_SIGNED(-501,11),
TO_SIGNED(-466,11),
TO_SIGNED(-428,11),
TO_SIGNED(-388,11),
TO_SIGNED(-347,11),
TO_SIGNED(-305,11),
TO_SIGNED(-262,11),
TO_SIGNED(-217,11),
TO_SIGNED(-172,11),
TO_SIGNED(-125,11),
TO_SIGNED(-79,11),
TO_SIGNED(-32,11),
TO_SIGNED(15,11),
TO_SIGNED(62,11),
TO_SIGNED(109,11),
TO_SIGNED(155,11),
TO_SIGNED(201,11),
TO_SIGNED(245,11),
TO_SIGNED(289,11),
TO_SIGNED(332,11),
TO_SIGNED(374,11),
TO_SIGNED(414,11),
TO_SIGNED(452,11),
TO_SIGNED(489,11),
TO_SIGNED(523,11),
TO_SIGNED(556,11),
TO_SIGNED(586,11),
TO_SIGNED(615,11),
TO_SIGNED(640,11),
TO_SIGNED(663,11),
TO_SIGNED(684,11),
TO_SIGNED(702,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(710,11),
TO_SIGNED(693,11),
TO_SIGNED(674,11),
TO_SIGNED(652,11),
TO_SIGNED(627,11),
TO_SIGNED(600,11),
TO_SIGNED(571,11),
TO_SIGNED(539,11),
TO_SIGNED(505,11),
TO_SIGNED(470,11),
TO_SIGNED(432,11),
TO_SIGNED(393,11),
TO_SIGNED(352,11),
TO_SIGNED(310,11),
TO_SIGNED(267,11),
TO_SIGNED(222,11),
TO_SIGNED(177,11),
TO_SIGNED(131,11),
TO_SIGNED(84,11),
TO_SIGNED(37,11),
TO_SIGNED(-10,11),
TO_SIGNED(-57,11),
TO_SIGNED(-103,11),
TO_SIGNED(-150,11),
TO_SIGNED(-195,11),
TO_SIGNED(-240,11),
TO_SIGNED(-284,11),
TO_SIGNED(-327,11),
TO_SIGNED(-369,11),
TO_SIGNED(-409,11),
TO_SIGNED(-448,11),
TO_SIGNED(-485,11),
TO_SIGNED(-519,11),
TO_SIGNED(-552,11),
TO_SIGNED(-583,11),
TO_SIGNED(-611,11),
TO_SIGNED(-637,11),
TO_SIGNED(-661,11),
TO_SIGNED(-682,11),
TO_SIGNED(-700,11),
TO_SIGNED(-716,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-725,11),
TO_SIGNED(-711,11),
TO_SIGNED(-695,11),
TO_SIGNED(-676,11),
TO_SIGNED(-654,11),
TO_SIGNED(-630,11),
TO_SIGNED(-603,11),
TO_SIGNED(-574,11),
TO_SIGNED(-543,11),
TO_SIGNED(-509,11),
TO_SIGNED(-474,11),
TO_SIGNED(-437,11),
TO_SIGNED(-397,11),
TO_SIGNED(-357,11),
TO_SIGNED(-315,11),
TO_SIGNED(-272,11),
TO_SIGNED(-227,11),
TO_SIGNED(-182,11),
TO_SIGNED(-136,11),
TO_SIGNED(-90,11),
TO_SIGNED(-43,11),
TO_SIGNED(4,11),
TO_SIGNED(51,11),
TO_SIGNED(98,11),
TO_SIGNED(144,11),
TO_SIGNED(190,11),
TO_SIGNED(235,11),
TO_SIGNED(279,11),
TO_SIGNED(323,11),
TO_SIGNED(364,11),
TO_SIGNED(405,11),
TO_SIGNED(443,11),
TO_SIGNED(480,11),
TO_SIGNED(516,11),
TO_SIGNED(549,11),
TO_SIGNED(580,11),
TO_SIGNED(608,11),
TO_SIGNED(635,11),
TO_SIGNED(658,11),
TO_SIGNED(680,11),
TO_SIGNED(698,11),
TO_SIGNED(714,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(713,11),
TO_SIGNED(697,11),
TO_SIGNED(678,11),
TO_SIGNED(657,11),
TO_SIGNED(633,11),
TO_SIGNED(606,11),
TO_SIGNED(578,11),
TO_SIGNED(547,11),
TO_SIGNED(513,11),
TO_SIGNED(478,11),
TO_SIGNED(441,11),
TO_SIGNED(402,11),
TO_SIGNED(362,11),
TO_SIGNED(320,11),
TO_SIGNED(276,11),
TO_SIGNED(232,11),
TO_SIGNED(187,11),
TO_SIGNED(141,11),
TO_SIGNED(95,11),
TO_SIGNED(48,11),
TO_SIGNED(1,11),
TO_SIGNED(-46,11),
TO_SIGNED(-93,11),
TO_SIGNED(-139,11),
TO_SIGNED(-185,11),
TO_SIGNED(-230,11),
TO_SIGNED(-275,11),
TO_SIGNED(-318,11),
TO_SIGNED(-360,11),
TO_SIGNED(-400,11),
TO_SIGNED(-439,11),
TO_SIGNED(-476,11),
TO_SIGNED(-512,11),
TO_SIGNED(-545,11),
TO_SIGNED(-576,11),
TO_SIGNED(-605,11),
TO_SIGNED(-632,11),
TO_SIGNED(-656,11),
TO_SIGNED(-677,11),
TO_SIGNED(-696,11),
TO_SIGNED(-712,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-715,11),
TO_SIGNED(-699,11),
TO_SIGNED(-681,11),
TO_SIGNED(-659,11),
TO_SIGNED(-636,11),
TO_SIGNED(-610,11),
TO_SIGNED(-581,11),
TO_SIGNED(-550,11),
TO_SIGNED(-517,11),
TO_SIGNED(-482,11),
TO_SIGNED(-445,11),
TO_SIGNED(-406,11),
TO_SIGNED(-366,11),
TO_SIGNED(-324,11),
TO_SIGNED(-281,11),
TO_SIGNED(-237,11),
TO_SIGNED(-192,11),
TO_SIGNED(-147,11),
TO_SIGNED(-100,11),
TO_SIGNED(-53,11),
TO_SIGNED(-6,11),
TO_SIGNED(41,11),
TO_SIGNED(87,11),
TO_SIGNED(134,11),
TO_SIGNED(180,11),
TO_SIGNED(225,11),
TO_SIGNED(270,11),
TO_SIGNED(313,11),
TO_SIGNED(355,11),
TO_SIGNED(396,11),
TO_SIGNED(435,11),
TO_SIGNED(472,11),
TO_SIGNED(508,11),
TO_SIGNED(541,11),
TO_SIGNED(573,11),
TO_SIGNED(602,11),
TO_SIGNED(629,11),
TO_SIGNED(653,11),
TO_SIGNED(675,11),
TO_SIGNED(694,11),
TO_SIGNED(711,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(729,11),
TO_SIGNED(716,11),
TO_SIGNED(701,11),
TO_SIGNED(683,11),
TO_SIGNED(662,11),
TO_SIGNED(639,11),
TO_SIGNED(613,11),
TO_SIGNED(584,11),
TO_SIGNED(554,11),
TO_SIGNED(521,11),
TO_SIGNED(486,11),
TO_SIGNED(449,11),
TO_SIGNED(411,11),
TO_SIGNED(371,11),
TO_SIGNED(329,11),
TO_SIGNED(286,11),
TO_SIGNED(242,11),
TO_SIGNED(197,11),
TO_SIGNED(152,11),
TO_SIGNED(105,11),
TO_SIGNED(59,11),
TO_SIGNED(12,11),
TO_SIGNED(-35,11),
TO_SIGNED(-82,11),
TO_SIGNED(-129,11),
TO_SIGNED(-175,11),
TO_SIGNED(-220,11),
TO_SIGNED(-265,11),
TO_SIGNED(-308,11),
TO_SIGNED(-350,11),
TO_SIGNED(-391,11),
TO_SIGNED(-430,11),
TO_SIGNED(-468,11),
TO_SIGNED(-504,11),
TO_SIGNED(-538,11),
TO_SIGNED(-569,11),
TO_SIGNED(-599,11),
TO_SIGNED(-626,11),
TO_SIGNED(-651,11),
TO_SIGNED(-673,11),
TO_SIGNED(-692,11),
TO_SIGNED(-709,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-685,11),
TO_SIGNED(-664,11),
TO_SIGNED(-641,11),
TO_SIGNED(-616,11),
TO_SIGNED(-588,11),
TO_SIGNED(-557,11),
TO_SIGNED(-525,11),
TO_SIGNED(-490,11),
TO_SIGNED(-454,11),
TO_SIGNED(-415,11),
TO_SIGNED(-375,11),
TO_SIGNED(-334,11),
TO_SIGNED(-291,11),
TO_SIGNED(-247,11),
TO_SIGNED(-203,11),
TO_SIGNED(-157,11),
TO_SIGNED(-111,11),
TO_SIGNED(-64,11),
TO_SIGNED(-17,11),
TO_SIGNED(30,11),
TO_SIGNED(77,11),
TO_SIGNED(123,11),
TO_SIGNED(169,11),
TO_SIGNED(215,11),
TO_SIGNED(260,11),
TO_SIGNED(303,11),
TO_SIGNED(345,11),
TO_SIGNED(387,11),
TO_SIGNED(426,11),
TO_SIGNED(464,11),
TO_SIGNED(500,11),
TO_SIGNED(534,11),
TO_SIGNED(566,11),
TO_SIGNED(596,11),
TO_SIGNED(623,11),
TO_SIGNED(648,11),
TO_SIGNED(670,11),
TO_SIGNED(690,11),
TO_SIGNED(707,11),
TO_SIGNED(721,11),
TO_SIGNED(733,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(705,11),
TO_SIGNED(687,11),
TO_SIGNED(667,11),
TO_SIGNED(644,11),
TO_SIGNED(619,11),
TO_SIGNED(591,11),
TO_SIGNED(561,11),
TO_SIGNED(529,11),
TO_SIGNED(494,11),
TO_SIGNED(458,11),
TO_SIGNED(420,11),
TO_SIGNED(380,11),
TO_SIGNED(339,11),
TO_SIGNED(296,11),
TO_SIGNED(252,11),
TO_SIGNED(208,11),
TO_SIGNED(162,11),
TO_SIGNED(116,11),
TO_SIGNED(69,11),
TO_SIGNED(22,11),
TO_SIGNED(-25,11),
TO_SIGNED(-71,11),
TO_SIGNED(-118,11),
TO_SIGNED(-164,11),
TO_SIGNED(-210,11),
TO_SIGNED(-255,11),
TO_SIGNED(-298,11),
TO_SIGNED(-341,11),
TO_SIGNED(-382,11),
TO_SIGNED(-422,11),
TO_SIGNED(-460,11),
TO_SIGNED(-496,11),
TO_SIGNED(-530,11),
TO_SIGNED(-562,11),
TO_SIGNED(-592,11),
TO_SIGNED(-620,11),
TO_SIGNED(-645,11),
TO_SIGNED(-668,11),
TO_SIGNED(-688,11),
TO_SIGNED(-705,11),
TO_SIGNED(-720,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-721,11),
TO_SIGNED(-706,11),
TO_SIGNED(-689,11),
TO_SIGNED(-669,11),
TO_SIGNED(-647,11),
TO_SIGNED(-622,11),
TO_SIGNED(-594,11),
TO_SIGNED(-564,11),
TO_SIGNED(-532,11),
TO_SIGNED(-498,11),
TO_SIGNED(-462,11),
TO_SIGNED(-424,11),
TO_SIGNED(-385,11),
TO_SIGNED(-344,11),
TO_SIGNED(-301,11),
TO_SIGNED(-258,11),
TO_SIGNED(-213,11),
TO_SIGNED(-167,11),
TO_SIGNED(-121,11),
TO_SIGNED(-75,11),
TO_SIGNED(-28,11),
TO_SIGNED(19,11),
TO_SIGNED(66,11),
TO_SIGNED(113,11),
TO_SIGNED(159,11),
TO_SIGNED(205,11),
TO_SIGNED(249,11),
TO_SIGNED(293,11),
TO_SIGNED(336,11),
TO_SIGNED(377,11),
TO_SIGNED(417,11),
TO_SIGNED(455,11),
TO_SIGNED(492,11),
TO_SIGNED(526,11),
TO_SIGNED(559,11),
TO_SIGNED(589,11),
TO_SIGNED(617,11),
TO_SIGNED(642,11),
TO_SIGNED(665,11),
TO_SIGNED(686,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(708,11),
TO_SIGNED(691,11),
TO_SIGNED(672,11),
TO_SIGNED(650,11),
TO_SIGNED(625,11),
TO_SIGNED(598,11),
TO_SIGNED(568,11),
TO_SIGNED(536,11),
TO_SIGNED(502,11),
TO_SIGNED(466,11),
TO_SIGNED(429,11),
TO_SIGNED(389,11),
TO_SIGNED(348,11),
TO_SIGNED(306,11),
TO_SIGNED(263,11),
TO_SIGNED(218,11),
TO_SIGNED(173,11),
TO_SIGNED(127,11),
TO_SIGNED(80,11),
TO_SIGNED(33,11),
TO_SIGNED(-14,11),
TO_SIGNED(-61,11),
TO_SIGNED(-108,11),
TO_SIGNED(-154,11),
TO_SIGNED(-200,11),
TO_SIGNED(-244,11),
TO_SIGNED(-288,11),
TO_SIGNED(-331,11),
TO_SIGNED(-373,11),
TO_SIGNED(-413,11),
TO_SIGNED(-451,11),
TO_SIGNED(-488,11),
TO_SIGNED(-523,11),
TO_SIGNED(-555,11),
TO_SIGNED(-586,11),
TO_SIGNED(-614,11),
TO_SIGNED(-640,11),
TO_SIGNED(-663,11),
TO_SIGNED(-684,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-729,11),
TO_SIGNED(-739,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-710,11),
TO_SIGNED(-693,11),
TO_SIGNED(-674,11),
TO_SIGNED(-652,11),
TO_SIGNED(-628,11),
TO_SIGNED(-601,11),
TO_SIGNED(-571,11),
TO_SIGNED(-540,11),
TO_SIGNED(-506,11),
TO_SIGNED(-471,11),
TO_SIGNED(-433,11),
TO_SIGNED(-394,11),
TO_SIGNED(-353,11),
TO_SIGNED(-311,11),
TO_SIGNED(-268,11),
TO_SIGNED(-223,11),
TO_SIGNED(-178,11),
TO_SIGNED(-132,11),
TO_SIGNED(-85,11),
TO_SIGNED(-38,11),
TO_SIGNED(9,11),
TO_SIGNED(56,11),
TO_SIGNED(102,11),
TO_SIGNED(149,11),
TO_SIGNED(194,11),
TO_SIGNED(239,11),
TO_SIGNED(283,11),
TO_SIGNED(326,11),
TO_SIGNED(368,11),
TO_SIGNED(408,11),
TO_SIGNED(447,11),
TO_SIGNED(484,11),
TO_SIGNED(519,11),
TO_SIGNED(552,11),
TO_SIGNED(582,11),
TO_SIGNED(611,11),
TO_SIGNED(637,11),
TO_SIGNED(660,11),
TO_SIGNED(681,11),
TO_SIGNED(700,11),
TO_SIGNED(715,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(736,11),
TO_SIGNED(725,11),
TO_SIGNED(712,11),
TO_SIGNED(695,11),
TO_SIGNED(676,11),
TO_SIGNED(655,11),
TO_SIGNED(631,11),
TO_SIGNED(604,11),
TO_SIGNED(575,11),
TO_SIGNED(544,11),
TO_SIGNED(510,11),
TO_SIGNED(475,11),
TO_SIGNED(437,11),
TO_SIGNED(398,11),
TO_SIGNED(358,11),
TO_SIGNED(316,11),
TO_SIGNED(273,11),
TO_SIGNED(228,11),
TO_SIGNED(183,11),
TO_SIGNED(137,11),
TO_SIGNED(91,11),
TO_SIGNED(44,11),
TO_SIGNED(-3,11),
TO_SIGNED(-50,11),
TO_SIGNED(-97,11),
TO_SIGNED(-143,11),
TO_SIGNED(-189,11),
TO_SIGNED(-234,11),
TO_SIGNED(-278,11),
TO_SIGNED(-322,11),
TO_SIGNED(-363,11),
TO_SIGNED(-404,11),
TO_SIGNED(-443,11),
TO_SIGNED(-480,11),
TO_SIGNED(-515,11),
TO_SIGNED(-548,11),
TO_SIGNED(-579,11),
TO_SIGNED(-608,11),
TO_SIGNED(-634,11),
TO_SIGNED(-658,11),
TO_SIGNED(-679,11),
TO_SIGNED(-698,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-679,11),
TO_SIGNED(-657,11),
TO_SIGNED(-633,11),
TO_SIGNED(-607,11),
TO_SIGNED(-578,11),
TO_SIGNED(-547,11),
TO_SIGNED(-514,11),
TO_SIGNED(-479,11),
TO_SIGNED(-442,11),
TO_SIGNED(-403,11),
TO_SIGNED(-362,11),
TO_SIGNED(-321,11),
TO_SIGNED(-277,11),
TO_SIGNED(-233,11),
TO_SIGNED(-188,11),
TO_SIGNED(-142,11),
TO_SIGNED(-96,11),
TO_SIGNED(-49,11),
TO_SIGNED(-2,11),
TO_SIGNED(45,11),
TO_SIGNED(92,11),
TO_SIGNED(138,11),
TO_SIGNED(184,11),
TO_SIGNED(229,11),
TO_SIGNED(274,11),
TO_SIGNED(317,11),
TO_SIGNED(359,11),
TO_SIGNED(399,11),
TO_SIGNED(438,11),
TO_SIGNED(476,11),
TO_SIGNED(511,11),
TO_SIGNED(544,11),
TO_SIGNED(576,11),
TO_SIGNED(605,11),
TO_SIGNED(631,11),
TO_SIGNED(655,11),
TO_SIGNED(677,11),
TO_SIGNED(696,11),
TO_SIGNED(712,11),
TO_SIGNED(725,11),
TO_SIGNED(736,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(715,11),
TO_SIGNED(699,11),
TO_SIGNED(681,11),
TO_SIGNED(660,11),
TO_SIGNED(636,11),
TO_SIGNED(610,11),
TO_SIGNED(582,11),
TO_SIGNED(551,11),
TO_SIGNED(518,11),
TO_SIGNED(483,11),
TO_SIGNED(446,11),
TO_SIGNED(407,11),
TO_SIGNED(367,11),
TO_SIGNED(325,11),
TO_SIGNED(282,11),
TO_SIGNED(238,11),
TO_SIGNED(193,11),
TO_SIGNED(148,11),
TO_SIGNED(101,11),
TO_SIGNED(54,11),
TO_SIGNED(7,11),
TO_SIGNED(-40,11),
TO_SIGNED(-86,11),
TO_SIGNED(-133,11),
TO_SIGNED(-179,11),
TO_SIGNED(-224,11),
TO_SIGNED(-269,11),
TO_SIGNED(-312,11),
TO_SIGNED(-354,11),
TO_SIGNED(-395,11),
TO_SIGNED(-434,11),
TO_SIGNED(-471,11),
TO_SIGNED(-507,11),
TO_SIGNED(-541,11),
TO_SIGNED(-572,11),
TO_SIGNED(-601,11),
TO_SIGNED(-628,11),
TO_SIGNED(-653,11),
TO_SIGNED(-675,11),
TO_SIGNED(-694,11),
TO_SIGNED(-710,11),
TO_SIGNED(-724,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-701,11),
TO_SIGNED(-683,11),
TO_SIGNED(-662,11),
TO_SIGNED(-639,11),
TO_SIGNED(-613,11),
TO_SIGNED(-585,11),
TO_SIGNED(-554,11),
TO_SIGNED(-522,11),
TO_SIGNED(-487,11),
TO_SIGNED(-450,11),
TO_SIGNED(-412,11),
TO_SIGNED(-372,11),
TO_SIGNED(-330,11),
TO_SIGNED(-287,11),
TO_SIGNED(-243,11),
TO_SIGNED(-198,11),
TO_SIGNED(-153,11),
TO_SIGNED(-106,11),
TO_SIGNED(-60,11),
TO_SIGNED(-13,11),
TO_SIGNED(34,11),
TO_SIGNED(81,11),
TO_SIGNED(128,11),
TO_SIGNED(174,11),
TO_SIGNED(219,11),
TO_SIGNED(264,11),
TO_SIGNED(307,11),
TO_SIGNED(349,11),
TO_SIGNED(390,11),
TO_SIGNED(430,11),
TO_SIGNED(467,11),
TO_SIGNED(503,11),
TO_SIGNED(537,11),
TO_SIGNED(569,11),
TO_SIGNED(598,11),
TO_SIGNED(625,11),
TO_SIGNED(650,11),
TO_SIGNED(672,11),
TO_SIGNED(692,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(730,11),
TO_SIGNED(718,11),
TO_SIGNED(703,11),
TO_SIGNED(685,11),
TO_SIGNED(665,11),
TO_SIGNED(642,11),
TO_SIGNED(616,11),
TO_SIGNED(588,11),
TO_SIGNED(558,11),
TO_SIGNED(526,11),
TO_SIGNED(491,11),
TO_SIGNED(455,11),
TO_SIGNED(416,11),
TO_SIGNED(376,11),
TO_SIGNED(335,11),
TO_SIGNED(292,11),
TO_SIGNED(248,11),
TO_SIGNED(204,11),
TO_SIGNED(158,11),
TO_SIGNED(112,11),
TO_SIGNED(65,11),
TO_SIGNED(18,11),
TO_SIGNED(-29,11),
TO_SIGNED(-76,11),
TO_SIGNED(-122,11),
TO_SIGNED(-168,11),
TO_SIGNED(-214,11),
TO_SIGNED(-259,11),
TO_SIGNED(-302,11),
TO_SIGNED(-345,11),
TO_SIGNED(-386,11),
TO_SIGNED(-425,11),
TO_SIGNED(-463,11),
TO_SIGNED(-499,11),
TO_SIGNED(-533,11),
TO_SIGNED(-565,11),
TO_SIGNED(-595,11),
TO_SIGNED(-622,11),
TO_SIGNED(-647,11),
TO_SIGNED(-670,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-721,11),
TO_SIGNED(-733,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-720,11),
TO_SIGNED(-705,11),
TO_SIGNED(-688,11),
TO_SIGNED(-667,11),
TO_SIGNED(-645,11),
TO_SIGNED(-619,11),
TO_SIGNED(-592,11),
TO_SIGNED(-562,11),
TO_SIGNED(-529,11),
TO_SIGNED(-495,11),
TO_SIGNED(-459,11),
TO_SIGNED(-421,11),
TO_SIGNED(-381,11),
TO_SIGNED(-340,11),
TO_SIGNED(-297,11),
TO_SIGNED(-254,11),
TO_SIGNED(-209,11),
TO_SIGNED(-163,11),
TO_SIGNED(-117,11),
TO_SIGNED(-70,11),
TO_SIGNED(-24,11),
TO_SIGNED(24,11),
TO_SIGNED(70,11),
TO_SIGNED(117,11),
TO_SIGNED(163,11),
TO_SIGNED(209,11),
TO_SIGNED(254,11),
TO_SIGNED(297,11),
TO_SIGNED(340,11),
TO_SIGNED(381,11),
TO_SIGNED(421,11),
TO_SIGNED(459,11),
TO_SIGNED(495,11),
TO_SIGNED(529,11),
TO_SIGNED(562,11),
TO_SIGNED(592,11),
TO_SIGNED(619,11),
TO_SIGNED(645,11),
TO_SIGNED(667,11),
TO_SIGNED(688,11),
TO_SIGNED(705,11),
TO_SIGNED(720,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(733,11),
TO_SIGNED(721,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(670,11),
TO_SIGNED(647,11),
TO_SIGNED(622,11),
TO_SIGNED(595,11),
TO_SIGNED(565,11),
TO_SIGNED(533,11),
TO_SIGNED(499,11),
TO_SIGNED(463,11),
TO_SIGNED(425,11),
TO_SIGNED(386,11),
TO_SIGNED(345,11),
TO_SIGNED(302,11),
TO_SIGNED(259,11),
TO_SIGNED(214,11),
TO_SIGNED(168,11),
TO_SIGNED(122,11),
TO_SIGNED(76,11),
TO_SIGNED(29,11),
TO_SIGNED(-18,11),
TO_SIGNED(-65,11),
TO_SIGNED(-112,11),
TO_SIGNED(-158,11),
TO_SIGNED(-204,11),
TO_SIGNED(-248,11),
TO_SIGNED(-292,11),
TO_SIGNED(-335,11),
TO_SIGNED(-376,11),
TO_SIGNED(-416,11),
TO_SIGNED(-455,11),
TO_SIGNED(-491,11),
TO_SIGNED(-526,11),
TO_SIGNED(-558,11),
TO_SIGNED(-588,11),
TO_SIGNED(-616,11),
TO_SIGNED(-642,11),
TO_SIGNED(-665,11),
TO_SIGNED(-685,11),
TO_SIGNED(-703,11),
TO_SIGNED(-718,11),
TO_SIGNED(-730,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-692,11),
TO_SIGNED(-672,11),
TO_SIGNED(-650,11),
TO_SIGNED(-625,11),
TO_SIGNED(-598,11),
TO_SIGNED(-569,11),
TO_SIGNED(-537,11),
TO_SIGNED(-503,11),
TO_SIGNED(-467,11),
TO_SIGNED(-430,11),
TO_SIGNED(-390,11),
TO_SIGNED(-349,11),
TO_SIGNED(-307,11),
TO_SIGNED(-264,11),
TO_SIGNED(-219,11),
TO_SIGNED(-174,11),
TO_SIGNED(-128,11),
TO_SIGNED(-81,11),
TO_SIGNED(-34,11),
TO_SIGNED(13,11),
TO_SIGNED(60,11),
TO_SIGNED(106,11),
TO_SIGNED(153,11),
TO_SIGNED(198,11),
TO_SIGNED(243,11),
TO_SIGNED(287,11),
TO_SIGNED(330,11),
TO_SIGNED(372,11),
TO_SIGNED(412,11),
TO_SIGNED(450,11),
TO_SIGNED(487,11),
TO_SIGNED(522,11),
TO_SIGNED(554,11),
TO_SIGNED(585,11),
TO_SIGNED(613,11),
TO_SIGNED(639,11),
TO_SIGNED(662,11),
TO_SIGNED(683,11),
TO_SIGNED(701,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(724,11),
TO_SIGNED(710,11),
TO_SIGNED(694,11),
TO_SIGNED(675,11),
TO_SIGNED(653,11),
TO_SIGNED(628,11),
TO_SIGNED(601,11),
TO_SIGNED(572,11),
TO_SIGNED(541,11),
TO_SIGNED(507,11),
TO_SIGNED(471,11),
TO_SIGNED(434,11),
TO_SIGNED(395,11),
TO_SIGNED(354,11),
TO_SIGNED(312,11),
TO_SIGNED(269,11),
TO_SIGNED(224,11),
TO_SIGNED(179,11),
TO_SIGNED(133,11),
TO_SIGNED(86,11),
TO_SIGNED(40,11),
TO_SIGNED(-7,11),
TO_SIGNED(-54,11),
TO_SIGNED(-101,11),
TO_SIGNED(-148,11),
TO_SIGNED(-193,11),
TO_SIGNED(-238,11),
TO_SIGNED(-282,11),
TO_SIGNED(-325,11),
TO_SIGNED(-367,11),
TO_SIGNED(-407,11),
TO_SIGNED(-446,11),
TO_SIGNED(-483,11),
TO_SIGNED(-518,11),
TO_SIGNED(-551,11),
TO_SIGNED(-582,11),
TO_SIGNED(-610,11),
TO_SIGNED(-636,11),
TO_SIGNED(-660,11),
TO_SIGNED(-681,11),
TO_SIGNED(-699,11),
TO_SIGNED(-715,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-736,11),
TO_SIGNED(-725,11),
TO_SIGNED(-712,11),
TO_SIGNED(-696,11),
TO_SIGNED(-677,11),
TO_SIGNED(-655,11),
TO_SIGNED(-631,11),
TO_SIGNED(-605,11),
TO_SIGNED(-576,11),
TO_SIGNED(-544,11),
TO_SIGNED(-511,11),
TO_SIGNED(-476,11),
TO_SIGNED(-438,11),
TO_SIGNED(-399,11),
TO_SIGNED(-359,11),
TO_SIGNED(-317,11),
TO_SIGNED(-274,11),
TO_SIGNED(-229,11),
TO_SIGNED(-184,11),
TO_SIGNED(-138,11),
TO_SIGNED(-92,11),
TO_SIGNED(-45,11),
TO_SIGNED(2,11),
TO_SIGNED(49,11),
TO_SIGNED(96,11),
TO_SIGNED(142,11),
TO_SIGNED(188,11),
TO_SIGNED(233,11),
TO_SIGNED(277,11),
TO_SIGNED(321,11),
TO_SIGNED(362,11),
TO_SIGNED(403,11),
TO_SIGNED(442,11),
TO_SIGNED(479,11),
TO_SIGNED(514,11),
TO_SIGNED(547,11),
TO_SIGNED(578,11),
TO_SIGNED(607,11),
TO_SIGNED(633,11),
TO_SIGNED(657,11),
TO_SIGNED(679,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(698,11),
TO_SIGNED(679,11),
TO_SIGNED(658,11),
TO_SIGNED(634,11),
TO_SIGNED(608,11),
TO_SIGNED(579,11),
TO_SIGNED(548,11),
TO_SIGNED(515,11),
TO_SIGNED(480,11),
TO_SIGNED(443,11),
TO_SIGNED(404,11),
TO_SIGNED(363,11),
TO_SIGNED(322,11),
TO_SIGNED(278,11),
TO_SIGNED(234,11),
TO_SIGNED(189,11),
TO_SIGNED(143,11),
TO_SIGNED(97,11),
TO_SIGNED(50,11),
TO_SIGNED(3,11),
TO_SIGNED(-44,11),
TO_SIGNED(-91,11),
TO_SIGNED(-137,11),
TO_SIGNED(-183,11),
TO_SIGNED(-228,11),
TO_SIGNED(-273,11),
TO_SIGNED(-316,11),
TO_SIGNED(-358,11),
TO_SIGNED(-398,11),
TO_SIGNED(-437,11),
TO_SIGNED(-475,11),
TO_SIGNED(-510,11),
TO_SIGNED(-544,11),
TO_SIGNED(-575,11),
TO_SIGNED(-604,11),
TO_SIGNED(-631,11),
TO_SIGNED(-655,11),
TO_SIGNED(-676,11),
TO_SIGNED(-695,11),
TO_SIGNED(-712,11),
TO_SIGNED(-725,11),
TO_SIGNED(-736,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-715,11),
TO_SIGNED(-700,11),
TO_SIGNED(-681,11),
TO_SIGNED(-660,11),
TO_SIGNED(-637,11),
TO_SIGNED(-611,11),
TO_SIGNED(-582,11),
TO_SIGNED(-552,11),
TO_SIGNED(-519,11),
TO_SIGNED(-484,11),
TO_SIGNED(-447,11),
TO_SIGNED(-408,11),
TO_SIGNED(-368,11),
TO_SIGNED(-326,11),
TO_SIGNED(-283,11),
TO_SIGNED(-239,11),
TO_SIGNED(-194,11),
TO_SIGNED(-149,11),
TO_SIGNED(-102,11),
TO_SIGNED(-56,11),
TO_SIGNED(-9,11),
TO_SIGNED(38,11),
TO_SIGNED(85,11),
TO_SIGNED(132,11),
TO_SIGNED(178,11),
TO_SIGNED(223,11),
TO_SIGNED(268,11),
TO_SIGNED(311,11),
TO_SIGNED(353,11),
TO_SIGNED(394,11),
TO_SIGNED(433,11),
TO_SIGNED(471,11),
TO_SIGNED(506,11),
TO_SIGNED(540,11),
TO_SIGNED(571,11),
TO_SIGNED(601,11),
TO_SIGNED(628,11),
TO_SIGNED(652,11),
TO_SIGNED(674,11),
TO_SIGNED(693,11),
TO_SIGNED(710,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(739,11),
TO_SIGNED(729,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(684,11),
TO_SIGNED(663,11),
TO_SIGNED(640,11),
TO_SIGNED(614,11),
TO_SIGNED(586,11),
TO_SIGNED(555,11),
TO_SIGNED(523,11),
TO_SIGNED(488,11),
TO_SIGNED(451,11),
TO_SIGNED(413,11),
TO_SIGNED(373,11),
TO_SIGNED(331,11),
TO_SIGNED(288,11),
TO_SIGNED(244,11),
TO_SIGNED(200,11),
TO_SIGNED(154,11),
TO_SIGNED(108,11),
TO_SIGNED(61,11),
TO_SIGNED(14,11),
TO_SIGNED(-33,11),
TO_SIGNED(-80,11),
TO_SIGNED(-127,11),
TO_SIGNED(-173,11),
TO_SIGNED(-218,11),
TO_SIGNED(-263,11),
TO_SIGNED(-306,11),
TO_SIGNED(-348,11),
TO_SIGNED(-389,11),
TO_SIGNED(-429,11),
TO_SIGNED(-466,11),
TO_SIGNED(-502,11),
TO_SIGNED(-536,11),
TO_SIGNED(-568,11),
TO_SIGNED(-598,11),
TO_SIGNED(-625,11),
TO_SIGNED(-650,11),
TO_SIGNED(-672,11),
TO_SIGNED(-691,11),
TO_SIGNED(-708,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-686,11),
TO_SIGNED(-665,11),
TO_SIGNED(-642,11),
TO_SIGNED(-617,11),
TO_SIGNED(-589,11),
TO_SIGNED(-559,11),
TO_SIGNED(-526,11),
TO_SIGNED(-492,11),
TO_SIGNED(-455,11),
TO_SIGNED(-417,11),
TO_SIGNED(-377,11),
TO_SIGNED(-336,11),
TO_SIGNED(-293,11),
TO_SIGNED(-249,11),
TO_SIGNED(-205,11),
TO_SIGNED(-159,11),
TO_SIGNED(-113,11),
TO_SIGNED(-66,11),
TO_SIGNED(-19,11),
TO_SIGNED(28,11),
TO_SIGNED(75,11),
TO_SIGNED(121,11),
TO_SIGNED(167,11),
TO_SIGNED(213,11),
TO_SIGNED(258,11),
TO_SIGNED(301,11),
TO_SIGNED(344,11),
TO_SIGNED(385,11),
TO_SIGNED(424,11),
TO_SIGNED(462,11),
TO_SIGNED(498,11),
TO_SIGNED(532,11),
TO_SIGNED(564,11),
TO_SIGNED(594,11),
TO_SIGNED(622,11),
TO_SIGNED(647,11),
TO_SIGNED(669,11),
TO_SIGNED(689,11),
TO_SIGNED(706,11),
TO_SIGNED(721,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(720,11),
TO_SIGNED(705,11),
TO_SIGNED(688,11),
TO_SIGNED(668,11),
TO_SIGNED(645,11),
TO_SIGNED(620,11),
TO_SIGNED(592,11),
TO_SIGNED(562,11),
TO_SIGNED(530,11),
TO_SIGNED(496,11),
TO_SIGNED(460,11),
TO_SIGNED(422,11),
TO_SIGNED(382,11),
TO_SIGNED(341,11),
TO_SIGNED(298,11),
TO_SIGNED(255,11),
TO_SIGNED(210,11),
TO_SIGNED(164,11),
TO_SIGNED(118,11),
TO_SIGNED(71,11),
TO_SIGNED(25,11),
TO_SIGNED(-22,11),
TO_SIGNED(-69,11),
TO_SIGNED(-116,11),
TO_SIGNED(-162,11),
TO_SIGNED(-208,11),
TO_SIGNED(-252,11),
TO_SIGNED(-296,11),
TO_SIGNED(-339,11),
TO_SIGNED(-380,11),
TO_SIGNED(-420,11),
TO_SIGNED(-458,11),
TO_SIGNED(-494,11),
TO_SIGNED(-529,11),
TO_SIGNED(-561,11),
TO_SIGNED(-591,11),
TO_SIGNED(-619,11),
TO_SIGNED(-644,11),
TO_SIGNED(-667,11),
TO_SIGNED(-687,11),
TO_SIGNED(-705,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-733,11),
TO_SIGNED(-721,11),
TO_SIGNED(-707,11),
TO_SIGNED(-690,11),
TO_SIGNED(-670,11),
TO_SIGNED(-648,11),
TO_SIGNED(-623,11),
TO_SIGNED(-596,11),
TO_SIGNED(-566,11),
TO_SIGNED(-534,11),
TO_SIGNED(-500,11),
TO_SIGNED(-464,11),
TO_SIGNED(-426,11),
TO_SIGNED(-387,11),
TO_SIGNED(-345,11),
TO_SIGNED(-303,11),
TO_SIGNED(-260,11),
TO_SIGNED(-215,11),
TO_SIGNED(-169,11),
TO_SIGNED(-123,11),
TO_SIGNED(-77,11),
TO_SIGNED(-30,11),
TO_SIGNED(17,11),
TO_SIGNED(64,11),
TO_SIGNED(111,11),
TO_SIGNED(157,11),
TO_SIGNED(203,11),
TO_SIGNED(247,11),
TO_SIGNED(291,11),
TO_SIGNED(334,11),
TO_SIGNED(375,11),
TO_SIGNED(415,11),
TO_SIGNED(454,11),
TO_SIGNED(490,11),
TO_SIGNED(525,11),
TO_SIGNED(557,11),
TO_SIGNED(588,11),
TO_SIGNED(616,11),
TO_SIGNED(641,11),
TO_SIGNED(664,11),
TO_SIGNED(685,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(709,11),
TO_SIGNED(692,11),
TO_SIGNED(673,11),
TO_SIGNED(651,11),
TO_SIGNED(626,11),
TO_SIGNED(599,11),
TO_SIGNED(569,11),
TO_SIGNED(538,11),
TO_SIGNED(504,11),
TO_SIGNED(468,11),
TO_SIGNED(430,11),
TO_SIGNED(391,11),
TO_SIGNED(350,11),
TO_SIGNED(308,11),
TO_SIGNED(265,11),
TO_SIGNED(220,11),
TO_SIGNED(175,11),
TO_SIGNED(129,11),
TO_SIGNED(82,11),
TO_SIGNED(35,11),
TO_SIGNED(-12,11),
TO_SIGNED(-59,11),
TO_SIGNED(-105,11),
TO_SIGNED(-152,11),
TO_SIGNED(-197,11),
TO_SIGNED(-242,11),
TO_SIGNED(-286,11),
TO_SIGNED(-329,11),
TO_SIGNED(-371,11),
TO_SIGNED(-411,11),
TO_SIGNED(-449,11),
TO_SIGNED(-486,11),
TO_SIGNED(-521,11),
TO_SIGNED(-554,11),
TO_SIGNED(-584,11),
TO_SIGNED(-613,11),
TO_SIGNED(-639,11),
TO_SIGNED(-662,11),
TO_SIGNED(-683,11),
TO_SIGNED(-701,11),
TO_SIGNED(-716,11),
TO_SIGNED(-729,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-711,11),
TO_SIGNED(-694,11),
TO_SIGNED(-675,11),
TO_SIGNED(-653,11),
TO_SIGNED(-629,11),
TO_SIGNED(-602,11),
TO_SIGNED(-573,11),
TO_SIGNED(-541,11),
TO_SIGNED(-508,11),
TO_SIGNED(-472,11),
TO_SIGNED(-435,11),
TO_SIGNED(-396,11),
TO_SIGNED(-355,11),
TO_SIGNED(-313,11),
TO_SIGNED(-270,11),
TO_SIGNED(-225,11),
TO_SIGNED(-180,11),
TO_SIGNED(-134,11),
TO_SIGNED(-87,11),
TO_SIGNED(-41,11),
TO_SIGNED(6,11),
TO_SIGNED(53,11),
TO_SIGNED(100,11),
TO_SIGNED(147,11),
TO_SIGNED(192,11),
TO_SIGNED(237,11),
TO_SIGNED(281,11),
TO_SIGNED(324,11),
TO_SIGNED(366,11),
TO_SIGNED(406,11),
TO_SIGNED(445,11),
TO_SIGNED(482,11),
TO_SIGNED(517,11),
TO_SIGNED(550,11),
TO_SIGNED(581,11),
TO_SIGNED(610,11),
TO_SIGNED(636,11),
TO_SIGNED(659,11),
TO_SIGNED(681,11),
TO_SIGNED(699,11),
TO_SIGNED(715,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(712,11),
TO_SIGNED(696,11),
TO_SIGNED(677,11),
TO_SIGNED(656,11),
TO_SIGNED(632,11),
TO_SIGNED(605,11),
TO_SIGNED(576,11),
TO_SIGNED(545,11),
TO_SIGNED(512,11),
TO_SIGNED(476,11),
TO_SIGNED(439,11),
TO_SIGNED(400,11),
TO_SIGNED(360,11),
TO_SIGNED(318,11),
TO_SIGNED(275,11),
TO_SIGNED(230,11),
TO_SIGNED(185,11),
TO_SIGNED(139,11),
TO_SIGNED(93,11),
TO_SIGNED(46,11),
TO_SIGNED(-1,11),
TO_SIGNED(-48,11),
TO_SIGNED(-95,11),
TO_SIGNED(-141,11),
TO_SIGNED(-187,11),
TO_SIGNED(-232,11),
TO_SIGNED(-276,11),
TO_SIGNED(-320,11),
TO_SIGNED(-362,11),
TO_SIGNED(-402,11),
TO_SIGNED(-441,11),
TO_SIGNED(-478,11),
TO_SIGNED(-513,11),
TO_SIGNED(-547,11),
TO_SIGNED(-578,11),
TO_SIGNED(-606,11),
TO_SIGNED(-633,11),
TO_SIGNED(-657,11),
TO_SIGNED(-678,11),
TO_SIGNED(-697,11),
TO_SIGNED(-713,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-714,11),
TO_SIGNED(-698,11),
TO_SIGNED(-680,11),
TO_SIGNED(-658,11),
TO_SIGNED(-635,11),
TO_SIGNED(-608,11),
TO_SIGNED(-580,11),
TO_SIGNED(-549,11),
TO_SIGNED(-516,11),
TO_SIGNED(-480,11),
TO_SIGNED(-443,11),
TO_SIGNED(-405,11),
TO_SIGNED(-364,11),
TO_SIGNED(-323,11),
TO_SIGNED(-279,11),
TO_SIGNED(-235,11),
TO_SIGNED(-190,11),
TO_SIGNED(-144,11),
TO_SIGNED(-98,11),
TO_SIGNED(-51,11),
TO_SIGNED(-4,11),
TO_SIGNED(43,11),
TO_SIGNED(90,11),
TO_SIGNED(136,11),
TO_SIGNED(182,11),
TO_SIGNED(227,11),
TO_SIGNED(272,11),
TO_SIGNED(315,11),
TO_SIGNED(357,11),
TO_SIGNED(397,11),
TO_SIGNED(437,11),
TO_SIGNED(474,11),
TO_SIGNED(509,11),
TO_SIGNED(543,11),
TO_SIGNED(574,11),
TO_SIGNED(603,11),
TO_SIGNED(630,11),
TO_SIGNED(654,11),
TO_SIGNED(676,11),
TO_SIGNED(695,11),
TO_SIGNED(711,11),
TO_SIGNED(725,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(716,11),
TO_SIGNED(700,11),
TO_SIGNED(682,11),
TO_SIGNED(661,11),
TO_SIGNED(637,11),
TO_SIGNED(611,11),
TO_SIGNED(583,11),
TO_SIGNED(552,11),
TO_SIGNED(519,11),
TO_SIGNED(485,11),
TO_SIGNED(448,11),
TO_SIGNED(409,11),
TO_SIGNED(369,11),
TO_SIGNED(327,11),
TO_SIGNED(284,11),
TO_SIGNED(240,11),
TO_SIGNED(195,11),
TO_SIGNED(150,11),
TO_SIGNED(103,11),
TO_SIGNED(57,11),
TO_SIGNED(10,11),
TO_SIGNED(-37,11),
TO_SIGNED(-84,11),
TO_SIGNED(-131,11),
TO_SIGNED(-177,11),
TO_SIGNED(-222,11),
TO_SIGNED(-267,11),
TO_SIGNED(-310,11),
TO_SIGNED(-352,11),
TO_SIGNED(-393,11),
TO_SIGNED(-432,11),
TO_SIGNED(-470,11),
TO_SIGNED(-505,11),
TO_SIGNED(-539,11),
TO_SIGNED(-571,11),
TO_SIGNED(-600,11),
TO_SIGNED(-627,11),
TO_SIGNED(-652,11),
TO_SIGNED(-674,11),
TO_SIGNED(-693,11),
TO_SIGNED(-710,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-702,11),
TO_SIGNED(-684,11),
TO_SIGNED(-663,11),
TO_SIGNED(-640,11),
TO_SIGNED(-615,11),
TO_SIGNED(-586,11),
TO_SIGNED(-556,11),
TO_SIGNED(-523,11),
TO_SIGNED(-489,11),
TO_SIGNED(-452,11),
TO_SIGNED(-414,11),
TO_SIGNED(-374,11),
TO_SIGNED(-332,11),
TO_SIGNED(-289,11),
TO_SIGNED(-245,11),
TO_SIGNED(-201,11),
TO_SIGNED(-155,11),
TO_SIGNED(-109,11),
TO_SIGNED(-62,11),
TO_SIGNED(-15,11),
TO_SIGNED(32,11),
TO_SIGNED(79,11),
TO_SIGNED(125,11),
TO_SIGNED(172,11),
TO_SIGNED(217,11),
TO_SIGNED(262,11),
TO_SIGNED(305,11),
TO_SIGNED(347,11),
TO_SIGNED(388,11),
TO_SIGNED(428,11),
TO_SIGNED(466,11),
TO_SIGNED(501,11),
TO_SIGNED(535,11),
TO_SIGNED(567,11),
TO_SIGNED(597,11),
TO_SIGNED(624,11),
TO_SIGNED(649,11),
TO_SIGNED(671,11),
TO_SIGNED(691,11),
TO_SIGNED(708,11),
TO_SIGNED(722,11),
TO_SIGNED(733,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(704,11),
TO_SIGNED(686,11),
TO_SIGNED(666,11),
TO_SIGNED(643,11),
TO_SIGNED(618,11),
TO_SIGNED(590,11),
TO_SIGNED(559,11),
TO_SIGNED(527,11),
TO_SIGNED(493,11),
TO_SIGNED(456,11),
TO_SIGNED(418,11),
TO_SIGNED(378,11),
TO_SIGNED(337,11),
TO_SIGNED(294,11),
TO_SIGNED(250,11),
TO_SIGNED(206,11),
TO_SIGNED(160,11),
TO_SIGNED(114,11),
TO_SIGNED(67,11),
TO_SIGNED(20,11),
TO_SIGNED(-27,11),
TO_SIGNED(-74,11),
TO_SIGNED(-120,11),
TO_SIGNED(-166,11),
TO_SIGNED(-212,11),
TO_SIGNED(-257,11),
TO_SIGNED(-300,11),
TO_SIGNED(-343,11),
TO_SIGNED(-384,11),
TO_SIGNED(-423,11),
TO_SIGNED(-461,11),
TO_SIGNED(-497,11),
TO_SIGNED(-532,11),
TO_SIGNED(-564,11),
TO_SIGNED(-594,11),
TO_SIGNED(-621,11),
TO_SIGNED(-646,11),
TO_SIGNED(-669,11),
TO_SIGNED(-689,11),
TO_SIGNED(-706,11),
TO_SIGNED(-721,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-720,11),
TO_SIGNED(-706,11),
TO_SIGNED(-688,11),
TO_SIGNED(-668,11),
TO_SIGNED(-646,11),
TO_SIGNED(-621,11),
TO_SIGNED(-593,11),
TO_SIGNED(-563,11),
TO_SIGNED(-531,11),
TO_SIGNED(-497,11),
TO_SIGNED(-460,11),
TO_SIGNED(-422,11),
TO_SIGNED(-383,11),
TO_SIGNED(-342,11),
TO_SIGNED(-299,11),
TO_SIGNED(-256,11),
TO_SIGNED(-211,11),
TO_SIGNED(-165,11),
TO_SIGNED(-119,11),
TO_SIGNED(-73,11),
TO_SIGNED(-26,11),
TO_SIGNED(21,11),
TO_SIGNED(68,11),
TO_SIGNED(115,11),
TO_SIGNED(161,11),
TO_SIGNED(207,11),
TO_SIGNED(251,11),
TO_SIGNED(295,11),
TO_SIGNED(338,11),
TO_SIGNED(379,11),
TO_SIGNED(419,11),
TO_SIGNED(457,11),
TO_SIGNED(493,11),
TO_SIGNED(528,11),
TO_SIGNED(560,11),
TO_SIGNED(590,11),
TO_SIGNED(618,11),
TO_SIGNED(644,11),
TO_SIGNED(666,11),
TO_SIGNED(687,11),
TO_SIGNED(704,11),
TO_SIGNED(719,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(671,11),
TO_SIGNED(648,11),
TO_SIGNED(624,11),
TO_SIGNED(596,11),
TO_SIGNED(567,11),
TO_SIGNED(535,11),
TO_SIGNED(501,11),
TO_SIGNED(465,11),
TO_SIGNED(427,11),
TO_SIGNED(387,11),
TO_SIGNED(346,11),
TO_SIGNED(304,11),
TO_SIGNED(261,11),
TO_SIGNED(216,11),
TO_SIGNED(171,11),
TO_SIGNED(124,11),
TO_SIGNED(78,11),
TO_SIGNED(31,11),
TO_SIGNED(-16,11),
TO_SIGNED(-63,11),
TO_SIGNED(-110,11),
TO_SIGNED(-156,11),
TO_SIGNED(-202,11),
TO_SIGNED(-246,11),
TO_SIGNED(-290,11),
TO_SIGNED(-333,11),
TO_SIGNED(-375,11),
TO_SIGNED(-415,11),
TO_SIGNED(-453,11),
TO_SIGNED(-489,11),
TO_SIGNED(-524,11),
TO_SIGNED(-557,11),
TO_SIGNED(-587,11),
TO_SIGNED(-615,11),
TO_SIGNED(-641,11),
TO_SIGNED(-664,11),
TO_SIGNED(-685,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-730,11),
TO_SIGNED(-739,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-693,11),
TO_SIGNED(-673,11),
TO_SIGNED(-651,11),
TO_SIGNED(-627,11),
TO_SIGNED(-599,11),
TO_SIGNED(-570,11),
TO_SIGNED(-538,11),
TO_SIGNED(-505,11),
TO_SIGNED(-469,11),
TO_SIGNED(-431,11),
TO_SIGNED(-392,11),
TO_SIGNED(-351,11),
TO_SIGNED(-309,11),
TO_SIGNED(-266,11),
TO_SIGNED(-221,11),
TO_SIGNED(-176,11),
TO_SIGNED(-130,11),
TO_SIGNED(-83,11),
TO_SIGNED(-36,11),
TO_SIGNED(11,11),
TO_SIGNED(58,11),
TO_SIGNED(104,11),
TO_SIGNED(151,11),
TO_SIGNED(196,11),
TO_SIGNED(241,11),
TO_SIGNED(285,11),
TO_SIGNED(328,11),
TO_SIGNED(370,11),
TO_SIGNED(410,11),
TO_SIGNED(449,11),
TO_SIGNED(485,11),
TO_SIGNED(520,11),
TO_SIGNED(553,11),
TO_SIGNED(584,11),
TO_SIGNED(612,11),
TO_SIGNED(638,11),
TO_SIGNED(661,11),
TO_SIGNED(682,11),
TO_SIGNED(700,11),
TO_SIGNED(716,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(725,11),
TO_SIGNED(711,11),
TO_SIGNED(695,11),
TO_SIGNED(675,11),
TO_SIGNED(654,11),
TO_SIGNED(629,11),
TO_SIGNED(603,11),
TO_SIGNED(574,11),
TO_SIGNED(542,11),
TO_SIGNED(509,11),
TO_SIGNED(473,11),
TO_SIGNED(436,11),
TO_SIGNED(397,11),
TO_SIGNED(356,11),
TO_SIGNED(314,11),
TO_SIGNED(271,11),
TO_SIGNED(226,11),
TO_SIGNED(181,11),
TO_SIGNED(135,11),
TO_SIGNED(88,11),
TO_SIGNED(42,11),
TO_SIGNED(-5,11),
TO_SIGNED(-52,11),
TO_SIGNED(-99,11),
TO_SIGNED(-145,11),
TO_SIGNED(-191,11),
TO_SIGNED(-236,11),
TO_SIGNED(-280,11),
TO_SIGNED(-323,11),
TO_SIGNED(-365,11),
TO_SIGNED(-406,11),
TO_SIGNED(-444,11),
TO_SIGNED(-481,11),
TO_SIGNED(-516,11),
TO_SIGNED(-549,11),
TO_SIGNED(-580,11),
TO_SIGNED(-609,11),
TO_SIGNED(-635,11),
TO_SIGNED(-659,11),
TO_SIGNED(-680,11),
TO_SIGNED(-699,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-736,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-678,11),
TO_SIGNED(-656,11),
TO_SIGNED(-632,11),
TO_SIGNED(-606,11),
TO_SIGNED(-577,11),
TO_SIGNED(-546,11),
TO_SIGNED(-512,11),
TO_SIGNED(-477,11),
TO_SIGNED(-440,11),
TO_SIGNED(-401,11),
TO_SIGNED(-361,11),
TO_SIGNED(-319,11),
TO_SIGNED(-275,11),
TO_SIGNED(-231,11),
TO_SIGNED(-186,11),
TO_SIGNED(-140,11),
TO_SIGNED(-94,11),
TO_SIGNED(-47,11),
TO_SIGNED(0,11),
TO_SIGNED(47,11),
TO_SIGNED(94,11),
TO_SIGNED(140,11),
TO_SIGNED(186,11),
TO_SIGNED(231,11),
TO_SIGNED(275,11),
TO_SIGNED(319,11),
TO_SIGNED(361,11),
TO_SIGNED(401,11),
TO_SIGNED(440,11),
TO_SIGNED(477,11),
TO_SIGNED(512,11),
TO_SIGNED(546,11),
TO_SIGNED(577,11),
TO_SIGNED(606,11),
TO_SIGNED(632,11),
TO_SIGNED(656,11),
TO_SIGNED(678,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(736,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(699,11),
TO_SIGNED(680,11),
TO_SIGNED(659,11),
TO_SIGNED(635,11),
TO_SIGNED(609,11),
TO_SIGNED(580,11),
TO_SIGNED(549,11),
TO_SIGNED(516,11),
TO_SIGNED(481,11),
TO_SIGNED(444,11),
TO_SIGNED(406,11),
TO_SIGNED(365,11),
TO_SIGNED(323,11),
TO_SIGNED(280,11),
TO_SIGNED(236,11),
TO_SIGNED(191,11),
TO_SIGNED(145,11),
TO_SIGNED(99,11),
TO_SIGNED(52,11),
TO_SIGNED(5,11),
TO_SIGNED(-42,11),
TO_SIGNED(-88,11),
TO_SIGNED(-135,11),
TO_SIGNED(-181,11),
TO_SIGNED(-226,11),
TO_SIGNED(-271,11),
TO_SIGNED(-314,11),
TO_SIGNED(-356,11),
TO_SIGNED(-397,11),
TO_SIGNED(-436,11),
TO_SIGNED(-473,11),
TO_SIGNED(-509,11),
TO_SIGNED(-542,11),
TO_SIGNED(-574,11),
TO_SIGNED(-603,11),
TO_SIGNED(-629,11),
TO_SIGNED(-654,11),
TO_SIGNED(-675,11),
TO_SIGNED(-695,11),
TO_SIGNED(-711,11),
TO_SIGNED(-725,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-716,11),
TO_SIGNED(-700,11),
TO_SIGNED(-682,11),
TO_SIGNED(-661,11),
TO_SIGNED(-638,11),
TO_SIGNED(-612,11),
TO_SIGNED(-584,11),
TO_SIGNED(-553,11),
TO_SIGNED(-520,11),
TO_SIGNED(-485,11),
TO_SIGNED(-449,11),
TO_SIGNED(-410,11),
TO_SIGNED(-370,11),
TO_SIGNED(-328,11),
TO_SIGNED(-285,11),
TO_SIGNED(-241,11),
TO_SIGNED(-196,11),
TO_SIGNED(-151,11),
TO_SIGNED(-104,11),
TO_SIGNED(-58,11),
TO_SIGNED(-11,11),
TO_SIGNED(36,11),
TO_SIGNED(83,11),
TO_SIGNED(130,11),
TO_SIGNED(176,11),
TO_SIGNED(221,11),
TO_SIGNED(266,11),
TO_SIGNED(309,11),
TO_SIGNED(351,11),
TO_SIGNED(392,11),
TO_SIGNED(431,11),
TO_SIGNED(469,11),
TO_SIGNED(505,11),
TO_SIGNED(538,11),
TO_SIGNED(570,11),
TO_SIGNED(599,11),
TO_SIGNED(627,11),
TO_SIGNED(651,11),
TO_SIGNED(673,11),
TO_SIGNED(693,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(739,11),
TO_SIGNED(730,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(685,11),
TO_SIGNED(664,11),
TO_SIGNED(641,11),
TO_SIGNED(615,11),
TO_SIGNED(587,11),
TO_SIGNED(557,11),
TO_SIGNED(524,11),
TO_SIGNED(489,11),
TO_SIGNED(453,11),
TO_SIGNED(415,11),
TO_SIGNED(375,11),
TO_SIGNED(333,11),
TO_SIGNED(290,11),
TO_SIGNED(246,11),
TO_SIGNED(202,11),
TO_SIGNED(156,11),
TO_SIGNED(110,11),
TO_SIGNED(63,11),
TO_SIGNED(16,11),
TO_SIGNED(-31,11),
TO_SIGNED(-78,11),
TO_SIGNED(-124,11),
TO_SIGNED(-171,11),
TO_SIGNED(-216,11),
TO_SIGNED(-261,11),
TO_SIGNED(-304,11),
TO_SIGNED(-346,11),
TO_SIGNED(-387,11),
TO_SIGNED(-427,11),
TO_SIGNED(-465,11),
TO_SIGNED(-501,11),
TO_SIGNED(-535,11),
TO_SIGNED(-567,11),
TO_SIGNED(-596,11),
TO_SIGNED(-624,11),
TO_SIGNED(-648,11),
TO_SIGNED(-671,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-719,11),
TO_SIGNED(-704,11),
TO_SIGNED(-687,11),
TO_SIGNED(-666,11),
TO_SIGNED(-644,11),
TO_SIGNED(-618,11),
TO_SIGNED(-590,11),
TO_SIGNED(-560,11),
TO_SIGNED(-528,11),
TO_SIGNED(-493,11),
TO_SIGNED(-457,11),
TO_SIGNED(-419,11),
TO_SIGNED(-379,11),
TO_SIGNED(-338,11),
TO_SIGNED(-295,11),
TO_SIGNED(-251,11),
TO_SIGNED(-207,11),
TO_SIGNED(-161,11),
TO_SIGNED(-115,11),
TO_SIGNED(-68,11),
TO_SIGNED(-21,11),
TO_SIGNED(26,11),
TO_SIGNED(73,11),
TO_SIGNED(119,11),
TO_SIGNED(165,11),
TO_SIGNED(211,11),
TO_SIGNED(256,11),
TO_SIGNED(299,11),
TO_SIGNED(342,11),
TO_SIGNED(383,11),
TO_SIGNED(422,11),
TO_SIGNED(460,11),
TO_SIGNED(497,11),
TO_SIGNED(531,11),
TO_SIGNED(563,11),
TO_SIGNED(593,11),
TO_SIGNED(621,11),
TO_SIGNED(646,11),
TO_SIGNED(668,11),
TO_SIGNED(688,11),
TO_SIGNED(706,11),
TO_SIGNED(720,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(721,11),
TO_SIGNED(706,11),
TO_SIGNED(689,11),
TO_SIGNED(669,11),
TO_SIGNED(646,11),
TO_SIGNED(621,11),
TO_SIGNED(594,11),
TO_SIGNED(564,11),
TO_SIGNED(532,11),
TO_SIGNED(497,11),
TO_SIGNED(461,11),
TO_SIGNED(423,11),
TO_SIGNED(384,11),
TO_SIGNED(343,11),
TO_SIGNED(300,11),
TO_SIGNED(257,11),
TO_SIGNED(212,11),
TO_SIGNED(166,11),
TO_SIGNED(120,11),
TO_SIGNED(74,11),
TO_SIGNED(27,11),
TO_SIGNED(-20,11),
TO_SIGNED(-67,11),
TO_SIGNED(-114,11),
TO_SIGNED(-160,11),
TO_SIGNED(-206,11),
TO_SIGNED(-250,11),
TO_SIGNED(-294,11),
TO_SIGNED(-337,11),
TO_SIGNED(-378,11),
TO_SIGNED(-418,11),
TO_SIGNED(-456,11),
TO_SIGNED(-493,11),
TO_SIGNED(-527,11),
TO_SIGNED(-559,11),
TO_SIGNED(-590,11),
TO_SIGNED(-618,11),
TO_SIGNED(-643,11),
TO_SIGNED(-666,11),
TO_SIGNED(-686,11),
TO_SIGNED(-704,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-733,11),
TO_SIGNED(-722,11),
TO_SIGNED(-708,11),
TO_SIGNED(-691,11),
TO_SIGNED(-671,11),
TO_SIGNED(-649,11),
TO_SIGNED(-624,11),
TO_SIGNED(-597,11),
TO_SIGNED(-567,11),
TO_SIGNED(-535,11),
TO_SIGNED(-501,11),
TO_SIGNED(-466,11),
TO_SIGNED(-428,11),
TO_SIGNED(-388,11),
TO_SIGNED(-347,11),
TO_SIGNED(-305,11),
TO_SIGNED(-262,11),
TO_SIGNED(-217,11),
TO_SIGNED(-172,11),
TO_SIGNED(-125,11),
TO_SIGNED(-79,11),
TO_SIGNED(-32,11),
TO_SIGNED(15,11),
TO_SIGNED(62,11),
TO_SIGNED(109,11),
TO_SIGNED(155,11),
TO_SIGNED(201,11),
TO_SIGNED(245,11),
TO_SIGNED(289,11),
TO_SIGNED(332,11),
TO_SIGNED(374,11),
TO_SIGNED(414,11),
TO_SIGNED(452,11),
TO_SIGNED(489,11),
TO_SIGNED(523,11),
TO_SIGNED(556,11),
TO_SIGNED(586,11),
TO_SIGNED(615,11),
TO_SIGNED(640,11),
TO_SIGNED(663,11),
TO_SIGNED(684,11),
TO_SIGNED(702,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(710,11),
TO_SIGNED(693,11),
TO_SIGNED(674,11),
TO_SIGNED(652,11),
TO_SIGNED(627,11),
TO_SIGNED(600,11),
TO_SIGNED(571,11),
TO_SIGNED(539,11),
TO_SIGNED(505,11),
TO_SIGNED(470,11),
TO_SIGNED(432,11),
TO_SIGNED(393,11),
TO_SIGNED(352,11),
TO_SIGNED(310,11),
TO_SIGNED(267,11),
TO_SIGNED(222,11),
TO_SIGNED(177,11),
TO_SIGNED(131,11),
TO_SIGNED(84,11),
TO_SIGNED(37,11),
TO_SIGNED(-10,11),
TO_SIGNED(-57,11),
TO_SIGNED(-103,11),
TO_SIGNED(-150,11),
TO_SIGNED(-195,11),
TO_SIGNED(-240,11),
TO_SIGNED(-284,11),
TO_SIGNED(-327,11),
TO_SIGNED(-369,11),
TO_SIGNED(-409,11),
TO_SIGNED(-448,11),
TO_SIGNED(-485,11),
TO_SIGNED(-519,11),
TO_SIGNED(-552,11),
TO_SIGNED(-583,11),
TO_SIGNED(-611,11),
TO_SIGNED(-637,11),
TO_SIGNED(-661,11),
TO_SIGNED(-682,11),
TO_SIGNED(-700,11),
TO_SIGNED(-716,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-725,11),
TO_SIGNED(-711,11),
TO_SIGNED(-695,11),
TO_SIGNED(-676,11),
TO_SIGNED(-654,11),
TO_SIGNED(-630,11),
TO_SIGNED(-603,11),
TO_SIGNED(-574,11),
TO_SIGNED(-543,11),
TO_SIGNED(-509,11),
TO_SIGNED(-474,11),
TO_SIGNED(-437,11),
TO_SIGNED(-397,11),
TO_SIGNED(-357,11),
TO_SIGNED(-315,11),
TO_SIGNED(-272,11),
TO_SIGNED(-227,11),
TO_SIGNED(-182,11),
TO_SIGNED(-136,11),
TO_SIGNED(-90,11),
TO_SIGNED(-43,11),
TO_SIGNED(4,11),
TO_SIGNED(51,11),
TO_SIGNED(98,11),
TO_SIGNED(144,11),
TO_SIGNED(190,11),
TO_SIGNED(235,11),
TO_SIGNED(279,11),
TO_SIGNED(323,11),
TO_SIGNED(364,11),
TO_SIGNED(405,11),
TO_SIGNED(443,11),
TO_SIGNED(480,11),
TO_SIGNED(516,11),
TO_SIGNED(549,11),
TO_SIGNED(580,11),
TO_SIGNED(608,11),
TO_SIGNED(635,11),
TO_SIGNED(658,11),
TO_SIGNED(680,11),
TO_SIGNED(698,11),
TO_SIGNED(714,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(713,11),
TO_SIGNED(697,11),
TO_SIGNED(678,11),
TO_SIGNED(657,11),
TO_SIGNED(633,11),
TO_SIGNED(606,11),
TO_SIGNED(578,11),
TO_SIGNED(547,11),
TO_SIGNED(513,11),
TO_SIGNED(478,11),
TO_SIGNED(441,11),
TO_SIGNED(402,11),
TO_SIGNED(362,11),
TO_SIGNED(320,11),
TO_SIGNED(276,11),
TO_SIGNED(232,11),
TO_SIGNED(187,11),
TO_SIGNED(141,11),
TO_SIGNED(95,11),
TO_SIGNED(48,11),
TO_SIGNED(1,11),
TO_SIGNED(-46,11),
TO_SIGNED(-93,11),
TO_SIGNED(-139,11),
TO_SIGNED(-185,11),
TO_SIGNED(-230,11),
TO_SIGNED(-275,11),
TO_SIGNED(-318,11),
TO_SIGNED(-360,11),
TO_SIGNED(-400,11),
TO_SIGNED(-439,11),
TO_SIGNED(-476,11),
TO_SIGNED(-512,11),
TO_SIGNED(-545,11),
TO_SIGNED(-576,11),
TO_SIGNED(-605,11),
TO_SIGNED(-632,11),
TO_SIGNED(-656,11),
TO_SIGNED(-677,11),
TO_SIGNED(-696,11),
TO_SIGNED(-712,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-715,11),
TO_SIGNED(-699,11),
TO_SIGNED(-681,11),
TO_SIGNED(-659,11),
TO_SIGNED(-636,11),
TO_SIGNED(-610,11),
TO_SIGNED(-581,11),
TO_SIGNED(-550,11),
TO_SIGNED(-517,11),
TO_SIGNED(-482,11),
TO_SIGNED(-445,11),
TO_SIGNED(-406,11),
TO_SIGNED(-366,11),
TO_SIGNED(-324,11),
TO_SIGNED(-281,11),
TO_SIGNED(-237,11),
TO_SIGNED(-192,11),
TO_SIGNED(-147,11),
TO_SIGNED(-100,11),
TO_SIGNED(-53,11),
TO_SIGNED(-6,11),
TO_SIGNED(41,11),
TO_SIGNED(87,11),
TO_SIGNED(134,11),
TO_SIGNED(180,11),
TO_SIGNED(225,11),
TO_SIGNED(270,11),
TO_SIGNED(313,11),
TO_SIGNED(355,11),
TO_SIGNED(396,11),
TO_SIGNED(435,11),
TO_SIGNED(472,11),
TO_SIGNED(508,11),
TO_SIGNED(541,11),
TO_SIGNED(573,11),
TO_SIGNED(602,11),
TO_SIGNED(629,11),
TO_SIGNED(653,11),
TO_SIGNED(675,11),
TO_SIGNED(694,11),
TO_SIGNED(711,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(729,11),
TO_SIGNED(716,11),
TO_SIGNED(701,11),
TO_SIGNED(683,11),
TO_SIGNED(662,11),
TO_SIGNED(639,11),
TO_SIGNED(613,11),
TO_SIGNED(584,11),
TO_SIGNED(554,11),
TO_SIGNED(521,11),
TO_SIGNED(486,11),
TO_SIGNED(449,11),
TO_SIGNED(411,11),
TO_SIGNED(371,11),
TO_SIGNED(329,11),
TO_SIGNED(286,11),
TO_SIGNED(242,11),
TO_SIGNED(197,11),
TO_SIGNED(152,11),
TO_SIGNED(105,11),
TO_SIGNED(59,11),
TO_SIGNED(12,11),
TO_SIGNED(-35,11),
TO_SIGNED(-82,11),
TO_SIGNED(-129,11),
TO_SIGNED(-175,11),
TO_SIGNED(-220,11),
TO_SIGNED(-265,11),
TO_SIGNED(-308,11),
TO_SIGNED(-350,11),
TO_SIGNED(-391,11),
TO_SIGNED(-430,11),
TO_SIGNED(-468,11),
TO_SIGNED(-504,11),
TO_SIGNED(-538,11),
TO_SIGNED(-569,11),
TO_SIGNED(-599,11),
TO_SIGNED(-626,11),
TO_SIGNED(-651,11),
TO_SIGNED(-673,11),
TO_SIGNED(-692,11),
TO_SIGNED(-709,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-685,11),
TO_SIGNED(-664,11),
TO_SIGNED(-641,11),
TO_SIGNED(-616,11),
TO_SIGNED(-588,11),
TO_SIGNED(-557,11),
TO_SIGNED(-525,11),
TO_SIGNED(-490,11),
TO_SIGNED(-454,11),
TO_SIGNED(-415,11),
TO_SIGNED(-375,11),
TO_SIGNED(-334,11),
TO_SIGNED(-291,11),
TO_SIGNED(-247,11),
TO_SIGNED(-203,11),
TO_SIGNED(-157,11),
TO_SIGNED(-111,11),
TO_SIGNED(-64,11),
TO_SIGNED(-17,11),
TO_SIGNED(30,11),
TO_SIGNED(77,11),
TO_SIGNED(123,11),
TO_SIGNED(169,11),
TO_SIGNED(215,11),
TO_SIGNED(260,11),
TO_SIGNED(303,11),
TO_SIGNED(345,11),
TO_SIGNED(387,11),
TO_SIGNED(426,11),
TO_SIGNED(464,11),
TO_SIGNED(500,11),
TO_SIGNED(534,11),
TO_SIGNED(566,11),
TO_SIGNED(596,11),
TO_SIGNED(623,11),
TO_SIGNED(648,11),
TO_SIGNED(670,11),
TO_SIGNED(690,11),
TO_SIGNED(707,11),
TO_SIGNED(721,11),
TO_SIGNED(733,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(705,11),
TO_SIGNED(687,11),
TO_SIGNED(667,11),
TO_SIGNED(644,11),
TO_SIGNED(619,11),
TO_SIGNED(591,11),
TO_SIGNED(561,11),
TO_SIGNED(529,11),
TO_SIGNED(494,11),
TO_SIGNED(458,11),
TO_SIGNED(420,11),
TO_SIGNED(380,11),
TO_SIGNED(339,11),
TO_SIGNED(296,11),
TO_SIGNED(252,11),
TO_SIGNED(208,11),
TO_SIGNED(162,11),
TO_SIGNED(116,11),
TO_SIGNED(69,11),
TO_SIGNED(22,11),
TO_SIGNED(-25,11),
TO_SIGNED(-71,11),
TO_SIGNED(-118,11),
TO_SIGNED(-164,11),
TO_SIGNED(-210,11),
TO_SIGNED(-255,11),
TO_SIGNED(-298,11),
TO_SIGNED(-341,11),
TO_SIGNED(-382,11),
TO_SIGNED(-422,11),
TO_SIGNED(-460,11),
TO_SIGNED(-496,11),
TO_SIGNED(-530,11),
TO_SIGNED(-562,11),
TO_SIGNED(-592,11),
TO_SIGNED(-620,11),
TO_SIGNED(-645,11),
TO_SIGNED(-668,11),
TO_SIGNED(-688,11),
TO_SIGNED(-705,11),
TO_SIGNED(-720,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-721,11),
TO_SIGNED(-706,11),
TO_SIGNED(-689,11),
TO_SIGNED(-669,11),
TO_SIGNED(-647,11),
TO_SIGNED(-622,11),
TO_SIGNED(-594,11),
TO_SIGNED(-564,11),
TO_SIGNED(-532,11),
TO_SIGNED(-498,11),
TO_SIGNED(-462,11),
TO_SIGNED(-424,11),
TO_SIGNED(-385,11),
TO_SIGNED(-344,11),
TO_SIGNED(-301,11),
TO_SIGNED(-258,11),
TO_SIGNED(-213,11),
TO_SIGNED(-167,11),
TO_SIGNED(-121,11),
TO_SIGNED(-75,11),
TO_SIGNED(-28,11),
TO_SIGNED(19,11),
TO_SIGNED(66,11),
TO_SIGNED(113,11),
TO_SIGNED(159,11),
TO_SIGNED(205,11),
TO_SIGNED(249,11),
TO_SIGNED(293,11),
TO_SIGNED(336,11),
TO_SIGNED(377,11),
TO_SIGNED(417,11),
TO_SIGNED(455,11),
TO_SIGNED(492,11),
TO_SIGNED(526,11),
TO_SIGNED(559,11),
TO_SIGNED(589,11),
TO_SIGNED(617,11),
TO_SIGNED(642,11),
TO_SIGNED(665,11),
TO_SIGNED(686,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(708,11),
TO_SIGNED(691,11),
TO_SIGNED(672,11),
TO_SIGNED(650,11),
TO_SIGNED(625,11),
TO_SIGNED(598,11),
TO_SIGNED(568,11),
TO_SIGNED(536,11),
TO_SIGNED(502,11),
TO_SIGNED(466,11),
TO_SIGNED(429,11),
TO_SIGNED(389,11),
TO_SIGNED(348,11),
TO_SIGNED(306,11),
TO_SIGNED(263,11),
TO_SIGNED(218,11),
TO_SIGNED(173,11),
TO_SIGNED(127,11),
TO_SIGNED(80,11),
TO_SIGNED(33,11),
TO_SIGNED(-14,11),
TO_SIGNED(-61,11),
TO_SIGNED(-108,11),
TO_SIGNED(-154,11),
TO_SIGNED(-200,11),
TO_SIGNED(-244,11),
TO_SIGNED(-288,11),
TO_SIGNED(-331,11),
TO_SIGNED(-373,11),
TO_SIGNED(-413,11),
TO_SIGNED(-451,11),
TO_SIGNED(-488,11),
TO_SIGNED(-523,11),
TO_SIGNED(-555,11),
TO_SIGNED(-586,11),
TO_SIGNED(-614,11),
TO_SIGNED(-640,11),
TO_SIGNED(-663,11),
TO_SIGNED(-684,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-729,11),
TO_SIGNED(-739,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-710,11),
TO_SIGNED(-693,11),
TO_SIGNED(-674,11),
TO_SIGNED(-652,11),
TO_SIGNED(-628,11),
TO_SIGNED(-601,11),
TO_SIGNED(-571,11),
TO_SIGNED(-540,11),
TO_SIGNED(-506,11),
TO_SIGNED(-471,11),
TO_SIGNED(-433,11),
TO_SIGNED(-394,11),
TO_SIGNED(-353,11),
TO_SIGNED(-311,11),
TO_SIGNED(-268,11),
TO_SIGNED(-223,11),
TO_SIGNED(-178,11),
TO_SIGNED(-132,11),
TO_SIGNED(-85,11),
TO_SIGNED(-38,11),
TO_SIGNED(9,11),
TO_SIGNED(56,11),
TO_SIGNED(102,11),
TO_SIGNED(149,11),
TO_SIGNED(194,11),
TO_SIGNED(239,11),
TO_SIGNED(283,11),
TO_SIGNED(326,11),
TO_SIGNED(368,11),
TO_SIGNED(408,11),
TO_SIGNED(447,11),
TO_SIGNED(484,11),
TO_SIGNED(519,11),
TO_SIGNED(552,11),
TO_SIGNED(582,11),
TO_SIGNED(611,11),
TO_SIGNED(637,11),
TO_SIGNED(660,11),
TO_SIGNED(681,11),
TO_SIGNED(700,11),
TO_SIGNED(715,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(736,11),
TO_SIGNED(725,11),
TO_SIGNED(712,11),
TO_SIGNED(695,11),
TO_SIGNED(676,11),
TO_SIGNED(655,11),
TO_SIGNED(631,11),
TO_SIGNED(604,11),
TO_SIGNED(575,11),
TO_SIGNED(544,11),
TO_SIGNED(510,11),
TO_SIGNED(475,11),
TO_SIGNED(437,11),
TO_SIGNED(398,11),
TO_SIGNED(358,11),
TO_SIGNED(316,11),
TO_SIGNED(273,11),
TO_SIGNED(228,11),
TO_SIGNED(183,11),
TO_SIGNED(137,11),
TO_SIGNED(91,11),
TO_SIGNED(44,11),
TO_SIGNED(-3,11),
TO_SIGNED(-50,11),
TO_SIGNED(-97,11),
TO_SIGNED(-143,11),
TO_SIGNED(-189,11),
TO_SIGNED(-234,11),
TO_SIGNED(-278,11),
TO_SIGNED(-322,11),
TO_SIGNED(-363,11),
TO_SIGNED(-404,11),
TO_SIGNED(-443,11),
TO_SIGNED(-480,11),
TO_SIGNED(-515,11),
TO_SIGNED(-548,11),
TO_SIGNED(-579,11),
TO_SIGNED(-608,11),
TO_SIGNED(-634,11),
TO_SIGNED(-658,11),
TO_SIGNED(-679,11),
TO_SIGNED(-698,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-679,11),
TO_SIGNED(-657,11),
TO_SIGNED(-633,11),
TO_SIGNED(-607,11),
TO_SIGNED(-578,11),
TO_SIGNED(-547,11),
TO_SIGNED(-514,11),
TO_SIGNED(-479,11),
TO_SIGNED(-442,11),
TO_SIGNED(-403,11),
TO_SIGNED(-362,11),
TO_SIGNED(-321,11),
TO_SIGNED(-277,11),
TO_SIGNED(-233,11),
TO_SIGNED(-188,11),
TO_SIGNED(-142,11),
TO_SIGNED(-96,11),
TO_SIGNED(-49,11),
TO_SIGNED(-2,11),
TO_SIGNED(45,11),
TO_SIGNED(92,11),
TO_SIGNED(138,11),
TO_SIGNED(184,11),
TO_SIGNED(229,11),
TO_SIGNED(274,11),
TO_SIGNED(317,11),
TO_SIGNED(359,11),
TO_SIGNED(399,11),
TO_SIGNED(438,11),
TO_SIGNED(476,11),
TO_SIGNED(511,11),
TO_SIGNED(544,11),
TO_SIGNED(576,11),
TO_SIGNED(605,11),
TO_SIGNED(631,11),
TO_SIGNED(655,11),
TO_SIGNED(677,11),
TO_SIGNED(696,11),
TO_SIGNED(712,11),
TO_SIGNED(725,11),
TO_SIGNED(736,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(715,11),
TO_SIGNED(699,11),
TO_SIGNED(681,11),
TO_SIGNED(660,11),
TO_SIGNED(636,11),
TO_SIGNED(610,11),
TO_SIGNED(582,11),
TO_SIGNED(551,11),
TO_SIGNED(518,11),
TO_SIGNED(483,11),
TO_SIGNED(446,11),
TO_SIGNED(407,11),
TO_SIGNED(367,11),
TO_SIGNED(325,11),
TO_SIGNED(282,11),
TO_SIGNED(238,11),
TO_SIGNED(193,11),
TO_SIGNED(148,11),
TO_SIGNED(101,11),
TO_SIGNED(54,11),
TO_SIGNED(7,11),
TO_SIGNED(-40,11),
TO_SIGNED(-86,11),
TO_SIGNED(-133,11),
TO_SIGNED(-179,11),
TO_SIGNED(-224,11),
TO_SIGNED(-269,11),
TO_SIGNED(-312,11),
TO_SIGNED(-354,11),
TO_SIGNED(-395,11),
TO_SIGNED(-434,11),
TO_SIGNED(-471,11),
TO_SIGNED(-507,11),
TO_SIGNED(-541,11),
TO_SIGNED(-572,11),
TO_SIGNED(-601,11),
TO_SIGNED(-628,11),
TO_SIGNED(-653,11),
TO_SIGNED(-675,11),
TO_SIGNED(-694,11),
TO_SIGNED(-710,11),
TO_SIGNED(-724,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-701,11),
TO_SIGNED(-683,11),
TO_SIGNED(-662,11),
TO_SIGNED(-639,11),
TO_SIGNED(-613,11),
TO_SIGNED(-585,11),
TO_SIGNED(-554,11),
TO_SIGNED(-522,11),
TO_SIGNED(-487,11),
TO_SIGNED(-450,11),
TO_SIGNED(-412,11),
TO_SIGNED(-372,11),
TO_SIGNED(-330,11),
TO_SIGNED(-287,11),
TO_SIGNED(-243,11),
TO_SIGNED(-198,11),
TO_SIGNED(-153,11),
TO_SIGNED(-106,11),
TO_SIGNED(-60,11),
TO_SIGNED(-13,11),
TO_SIGNED(34,11),
TO_SIGNED(81,11),
TO_SIGNED(128,11),
TO_SIGNED(174,11),
TO_SIGNED(219,11),
TO_SIGNED(264,11),
TO_SIGNED(307,11),
TO_SIGNED(349,11),
TO_SIGNED(390,11),
TO_SIGNED(430,11),
TO_SIGNED(467,11),
TO_SIGNED(503,11),
TO_SIGNED(537,11),
TO_SIGNED(569,11),
TO_SIGNED(598,11),
TO_SIGNED(625,11),
TO_SIGNED(650,11),
TO_SIGNED(672,11),
TO_SIGNED(692,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(730,11),
TO_SIGNED(718,11),
TO_SIGNED(703,11),
TO_SIGNED(685,11),
TO_SIGNED(665,11),
TO_SIGNED(642,11),
TO_SIGNED(616,11),
TO_SIGNED(588,11),
TO_SIGNED(558,11),
TO_SIGNED(526,11),
TO_SIGNED(491,11),
TO_SIGNED(455,11),
TO_SIGNED(416,11),
TO_SIGNED(376,11),
TO_SIGNED(335,11),
TO_SIGNED(292,11),
TO_SIGNED(248,11),
TO_SIGNED(204,11),
TO_SIGNED(158,11),
TO_SIGNED(112,11),
TO_SIGNED(65,11),
TO_SIGNED(18,11),
TO_SIGNED(-29,11),
TO_SIGNED(-76,11),
TO_SIGNED(-122,11),
TO_SIGNED(-168,11),
TO_SIGNED(-214,11),
TO_SIGNED(-259,11),
TO_SIGNED(-302,11),
TO_SIGNED(-345,11),
TO_SIGNED(-386,11),
TO_SIGNED(-425,11),
TO_SIGNED(-463,11),
TO_SIGNED(-499,11),
TO_SIGNED(-533,11),
TO_SIGNED(-565,11),
TO_SIGNED(-595,11),
TO_SIGNED(-622,11),
TO_SIGNED(-647,11),
TO_SIGNED(-670,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-721,11),
TO_SIGNED(-733,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-720,11),
TO_SIGNED(-705,11),
TO_SIGNED(-688,11),
TO_SIGNED(-667,11),
TO_SIGNED(-645,11),
TO_SIGNED(-619,11),
TO_SIGNED(-592,11),
TO_SIGNED(-562,11),
TO_SIGNED(-529,11),
TO_SIGNED(-495,11),
TO_SIGNED(-459,11),
TO_SIGNED(-421,11),
TO_SIGNED(-381,11),
TO_SIGNED(-340,11),
TO_SIGNED(-297,11),
TO_SIGNED(-254,11),
TO_SIGNED(-209,11),
TO_SIGNED(-163,11),
TO_SIGNED(-117,11),
TO_SIGNED(-70,11),
TO_SIGNED(-24,11),
TO_SIGNED(24,11),
TO_SIGNED(70,11),
TO_SIGNED(117,11),
TO_SIGNED(163,11),
TO_SIGNED(209,11),
TO_SIGNED(254,11),
TO_SIGNED(297,11),
TO_SIGNED(340,11),
TO_SIGNED(381,11),
TO_SIGNED(421,11),
TO_SIGNED(459,11),
TO_SIGNED(495,11),
TO_SIGNED(529,11),
TO_SIGNED(562,11),
TO_SIGNED(592,11),
TO_SIGNED(619,11),
TO_SIGNED(645,11),
TO_SIGNED(667,11),
TO_SIGNED(688,11),
TO_SIGNED(705,11),
TO_SIGNED(720,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(733,11),
TO_SIGNED(721,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(670,11),
TO_SIGNED(647,11),
TO_SIGNED(622,11),
TO_SIGNED(595,11),
TO_SIGNED(565,11),
TO_SIGNED(533,11),
TO_SIGNED(499,11),
TO_SIGNED(463,11),
TO_SIGNED(425,11),
TO_SIGNED(386,11),
TO_SIGNED(345,11),
TO_SIGNED(302,11),
TO_SIGNED(259,11),
TO_SIGNED(214,11),
TO_SIGNED(168,11),
TO_SIGNED(122,11),
TO_SIGNED(76,11),
TO_SIGNED(29,11),
TO_SIGNED(-18,11),
TO_SIGNED(-65,11),
TO_SIGNED(-112,11),
TO_SIGNED(-158,11),
TO_SIGNED(-204,11),
TO_SIGNED(-248,11),
TO_SIGNED(-292,11),
TO_SIGNED(-335,11),
TO_SIGNED(-376,11),
TO_SIGNED(-416,11),
TO_SIGNED(-455,11),
TO_SIGNED(-491,11),
TO_SIGNED(-526,11),
TO_SIGNED(-558,11),
TO_SIGNED(-588,11),
TO_SIGNED(-616,11),
TO_SIGNED(-642,11),
TO_SIGNED(-665,11),
TO_SIGNED(-685,11),
TO_SIGNED(-703,11),
TO_SIGNED(-718,11),
TO_SIGNED(-730,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-692,11),
TO_SIGNED(-672,11),
TO_SIGNED(-650,11),
TO_SIGNED(-625,11),
TO_SIGNED(-598,11),
TO_SIGNED(-569,11),
TO_SIGNED(-537,11),
TO_SIGNED(-503,11),
TO_SIGNED(-467,11),
TO_SIGNED(-430,11),
TO_SIGNED(-390,11),
TO_SIGNED(-349,11),
TO_SIGNED(-307,11),
TO_SIGNED(-264,11),
TO_SIGNED(-219,11),
TO_SIGNED(-174,11),
TO_SIGNED(-128,11),
TO_SIGNED(-81,11),
TO_SIGNED(-34,11),
TO_SIGNED(13,11),
TO_SIGNED(60,11),
TO_SIGNED(106,11),
TO_SIGNED(153,11),
TO_SIGNED(198,11),
TO_SIGNED(243,11),
TO_SIGNED(287,11),
TO_SIGNED(330,11),
TO_SIGNED(372,11),
TO_SIGNED(412,11),
TO_SIGNED(450,11),
TO_SIGNED(487,11),
TO_SIGNED(522,11),
TO_SIGNED(554,11),
TO_SIGNED(585,11),
TO_SIGNED(613,11),
TO_SIGNED(639,11),
TO_SIGNED(662,11),
TO_SIGNED(683,11),
TO_SIGNED(701,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(724,11),
TO_SIGNED(710,11),
TO_SIGNED(694,11),
TO_SIGNED(675,11),
TO_SIGNED(653,11),
TO_SIGNED(628,11),
TO_SIGNED(601,11),
TO_SIGNED(572,11),
TO_SIGNED(541,11),
TO_SIGNED(507,11),
TO_SIGNED(471,11),
TO_SIGNED(434,11),
TO_SIGNED(395,11),
TO_SIGNED(354,11),
TO_SIGNED(312,11),
TO_SIGNED(269,11),
TO_SIGNED(224,11),
TO_SIGNED(179,11),
TO_SIGNED(133,11),
TO_SIGNED(86,11),
TO_SIGNED(40,11),
TO_SIGNED(-7,11),
TO_SIGNED(-54,11),
TO_SIGNED(-101,11),
TO_SIGNED(-148,11),
TO_SIGNED(-193,11),
TO_SIGNED(-238,11),
TO_SIGNED(-282,11),
TO_SIGNED(-325,11),
TO_SIGNED(-367,11),
TO_SIGNED(-407,11),
TO_SIGNED(-446,11),
TO_SIGNED(-483,11),
TO_SIGNED(-518,11),
TO_SIGNED(-551,11),
TO_SIGNED(-582,11),
TO_SIGNED(-610,11),
TO_SIGNED(-636,11),
TO_SIGNED(-660,11),
TO_SIGNED(-681,11),
TO_SIGNED(-699,11),
TO_SIGNED(-715,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-736,11),
TO_SIGNED(-725,11),
TO_SIGNED(-712,11),
TO_SIGNED(-696,11),
TO_SIGNED(-677,11),
TO_SIGNED(-655,11),
TO_SIGNED(-631,11),
TO_SIGNED(-605,11),
TO_SIGNED(-576,11),
TO_SIGNED(-544,11),
TO_SIGNED(-511,11),
TO_SIGNED(-476,11),
TO_SIGNED(-438,11),
TO_SIGNED(-399,11),
TO_SIGNED(-359,11),
TO_SIGNED(-317,11),
TO_SIGNED(-274,11),
TO_SIGNED(-229,11),
TO_SIGNED(-184,11),
TO_SIGNED(-138,11),
TO_SIGNED(-92,11),
TO_SIGNED(-45,11),
TO_SIGNED(2,11),
TO_SIGNED(49,11),
TO_SIGNED(96,11),
TO_SIGNED(142,11),
TO_SIGNED(188,11),
TO_SIGNED(233,11),
TO_SIGNED(277,11),
TO_SIGNED(321,11),
TO_SIGNED(362,11),
TO_SIGNED(403,11),
TO_SIGNED(442,11),
TO_SIGNED(479,11),
TO_SIGNED(514,11),
TO_SIGNED(547,11),
TO_SIGNED(578,11),
TO_SIGNED(607,11),
TO_SIGNED(633,11),
TO_SIGNED(657,11),
TO_SIGNED(679,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(698,11),
TO_SIGNED(679,11),
TO_SIGNED(658,11),
TO_SIGNED(634,11),
TO_SIGNED(608,11),
TO_SIGNED(579,11),
TO_SIGNED(548,11),
TO_SIGNED(515,11),
TO_SIGNED(480,11),
TO_SIGNED(443,11),
TO_SIGNED(404,11),
TO_SIGNED(363,11),
TO_SIGNED(322,11),
TO_SIGNED(278,11),
TO_SIGNED(234,11),
TO_SIGNED(189,11),
TO_SIGNED(143,11),
TO_SIGNED(97,11),
TO_SIGNED(50,11),
TO_SIGNED(3,11),
TO_SIGNED(-44,11),
TO_SIGNED(-91,11),
TO_SIGNED(-137,11),
TO_SIGNED(-183,11),
TO_SIGNED(-228,11),
TO_SIGNED(-273,11),
TO_SIGNED(-316,11),
TO_SIGNED(-358,11),
TO_SIGNED(-398,11),
TO_SIGNED(-437,11),
TO_SIGNED(-475,11),
TO_SIGNED(-510,11),
TO_SIGNED(-544,11),
TO_SIGNED(-575,11),
TO_SIGNED(-604,11),
TO_SIGNED(-631,11),
TO_SIGNED(-655,11),
TO_SIGNED(-676,11),
TO_SIGNED(-695,11),
TO_SIGNED(-712,11),
TO_SIGNED(-725,11),
TO_SIGNED(-736,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-715,11),
TO_SIGNED(-700,11),
TO_SIGNED(-681,11),
TO_SIGNED(-660,11),
TO_SIGNED(-637,11),
TO_SIGNED(-611,11),
TO_SIGNED(-582,11),
TO_SIGNED(-552,11),
TO_SIGNED(-519,11),
TO_SIGNED(-484,11),
TO_SIGNED(-447,11),
TO_SIGNED(-408,11),
TO_SIGNED(-368,11),
TO_SIGNED(-326,11),
TO_SIGNED(-283,11),
TO_SIGNED(-239,11),
TO_SIGNED(-194,11),
TO_SIGNED(-149,11),
TO_SIGNED(-102,11),
TO_SIGNED(-56,11),
TO_SIGNED(-9,11),
TO_SIGNED(38,11),
TO_SIGNED(85,11),
TO_SIGNED(132,11),
TO_SIGNED(178,11),
TO_SIGNED(223,11),
TO_SIGNED(268,11),
TO_SIGNED(311,11),
TO_SIGNED(353,11),
TO_SIGNED(394,11),
TO_SIGNED(433,11),
TO_SIGNED(471,11),
TO_SIGNED(506,11),
TO_SIGNED(540,11),
TO_SIGNED(571,11),
TO_SIGNED(601,11),
TO_SIGNED(628,11),
TO_SIGNED(652,11),
TO_SIGNED(674,11),
TO_SIGNED(693,11),
TO_SIGNED(710,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(739,11),
TO_SIGNED(729,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(684,11),
TO_SIGNED(663,11),
TO_SIGNED(640,11),
TO_SIGNED(614,11),
TO_SIGNED(586,11),
TO_SIGNED(555,11),
TO_SIGNED(523,11),
TO_SIGNED(488,11),
TO_SIGNED(451,11),
TO_SIGNED(413,11),
TO_SIGNED(373,11),
TO_SIGNED(331,11),
TO_SIGNED(288,11),
TO_SIGNED(244,11),
TO_SIGNED(200,11),
TO_SIGNED(154,11),
TO_SIGNED(108,11),
TO_SIGNED(61,11),
TO_SIGNED(14,11),
TO_SIGNED(-33,11),
TO_SIGNED(-80,11),
TO_SIGNED(-127,11),
TO_SIGNED(-173,11),
TO_SIGNED(-218,11),
TO_SIGNED(-263,11),
TO_SIGNED(-306,11),
TO_SIGNED(-348,11),
TO_SIGNED(-389,11),
TO_SIGNED(-429,11),
TO_SIGNED(-466,11),
TO_SIGNED(-502,11),
TO_SIGNED(-536,11),
TO_SIGNED(-568,11),
TO_SIGNED(-598,11),
TO_SIGNED(-625,11),
TO_SIGNED(-650,11),
TO_SIGNED(-672,11),
TO_SIGNED(-691,11),
TO_SIGNED(-708,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-686,11),
TO_SIGNED(-665,11),
TO_SIGNED(-642,11),
TO_SIGNED(-617,11),
TO_SIGNED(-589,11),
TO_SIGNED(-559,11),
TO_SIGNED(-526,11),
TO_SIGNED(-492,11),
TO_SIGNED(-455,11),
TO_SIGNED(-417,11),
TO_SIGNED(-377,11),
TO_SIGNED(-336,11),
TO_SIGNED(-293,11),
TO_SIGNED(-249,11),
TO_SIGNED(-205,11),
TO_SIGNED(-159,11),
TO_SIGNED(-113,11),
TO_SIGNED(-66,11),
TO_SIGNED(-19,11),
TO_SIGNED(28,11),
TO_SIGNED(75,11),
TO_SIGNED(121,11),
TO_SIGNED(167,11),
TO_SIGNED(213,11),
TO_SIGNED(258,11),
TO_SIGNED(301,11),
TO_SIGNED(344,11),
TO_SIGNED(385,11),
TO_SIGNED(424,11),
TO_SIGNED(462,11),
TO_SIGNED(498,11),
TO_SIGNED(532,11),
TO_SIGNED(564,11),
TO_SIGNED(594,11),
TO_SIGNED(622,11),
TO_SIGNED(647,11),
TO_SIGNED(669,11),
TO_SIGNED(689,11),
TO_SIGNED(706,11),
TO_SIGNED(721,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(720,11),
TO_SIGNED(705,11),
TO_SIGNED(688,11),
TO_SIGNED(668,11),
TO_SIGNED(645,11),
TO_SIGNED(620,11),
TO_SIGNED(592,11),
TO_SIGNED(562,11),
TO_SIGNED(530,11),
TO_SIGNED(496,11),
TO_SIGNED(460,11),
TO_SIGNED(422,11),
TO_SIGNED(382,11),
TO_SIGNED(341,11),
TO_SIGNED(298,11),
TO_SIGNED(255,11),
TO_SIGNED(210,11),
TO_SIGNED(164,11),
TO_SIGNED(118,11),
TO_SIGNED(71,11),
TO_SIGNED(25,11),
TO_SIGNED(-22,11),
TO_SIGNED(-69,11),
TO_SIGNED(-116,11),
TO_SIGNED(-162,11),
TO_SIGNED(-208,11),
TO_SIGNED(-252,11),
TO_SIGNED(-296,11),
TO_SIGNED(-339,11),
TO_SIGNED(-380,11),
TO_SIGNED(-420,11),
TO_SIGNED(-458,11),
TO_SIGNED(-494,11),
TO_SIGNED(-529,11),
TO_SIGNED(-561,11),
TO_SIGNED(-591,11),
TO_SIGNED(-619,11),
TO_SIGNED(-644,11),
TO_SIGNED(-667,11),
TO_SIGNED(-687,11),
TO_SIGNED(-705,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-733,11),
TO_SIGNED(-721,11),
TO_SIGNED(-707,11),
TO_SIGNED(-690,11),
TO_SIGNED(-670,11),
TO_SIGNED(-648,11),
TO_SIGNED(-623,11),
TO_SIGNED(-596,11),
TO_SIGNED(-566,11),
TO_SIGNED(-534,11),
TO_SIGNED(-500,11),
TO_SIGNED(-464,11),
TO_SIGNED(-426,11),
TO_SIGNED(-387,11),
TO_SIGNED(-345,11),
TO_SIGNED(-303,11),
TO_SIGNED(-260,11),
TO_SIGNED(-215,11),
TO_SIGNED(-169,11),
TO_SIGNED(-123,11),
TO_SIGNED(-77,11),
TO_SIGNED(-30,11),
TO_SIGNED(17,11),
TO_SIGNED(64,11),
TO_SIGNED(111,11),
TO_SIGNED(157,11),
TO_SIGNED(203,11),
TO_SIGNED(247,11),
TO_SIGNED(291,11),
TO_SIGNED(334,11),
TO_SIGNED(375,11),
TO_SIGNED(415,11),
TO_SIGNED(454,11),
TO_SIGNED(490,11),
TO_SIGNED(525,11),
TO_SIGNED(557,11),
TO_SIGNED(588,11),
TO_SIGNED(616,11),
TO_SIGNED(641,11),
TO_SIGNED(664,11),
TO_SIGNED(685,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(709,11),
TO_SIGNED(692,11),
TO_SIGNED(673,11),
TO_SIGNED(651,11),
TO_SIGNED(626,11),
TO_SIGNED(599,11),
TO_SIGNED(569,11),
TO_SIGNED(538,11),
TO_SIGNED(504,11),
TO_SIGNED(468,11),
TO_SIGNED(430,11),
TO_SIGNED(391,11),
TO_SIGNED(350,11),
TO_SIGNED(308,11),
TO_SIGNED(265,11),
TO_SIGNED(220,11),
TO_SIGNED(175,11),
TO_SIGNED(129,11),
TO_SIGNED(82,11),
TO_SIGNED(35,11),
TO_SIGNED(-12,11),
TO_SIGNED(-59,11),
TO_SIGNED(-105,11),
TO_SIGNED(-152,11),
TO_SIGNED(-197,11),
TO_SIGNED(-242,11),
TO_SIGNED(-286,11),
TO_SIGNED(-329,11),
TO_SIGNED(-371,11),
TO_SIGNED(-411,11),
TO_SIGNED(-449,11),
TO_SIGNED(-486,11),
TO_SIGNED(-521,11),
TO_SIGNED(-554,11),
TO_SIGNED(-584,11),
TO_SIGNED(-613,11),
TO_SIGNED(-639,11),
TO_SIGNED(-662,11),
TO_SIGNED(-683,11),
TO_SIGNED(-701,11),
TO_SIGNED(-716,11),
TO_SIGNED(-729,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-711,11),
TO_SIGNED(-694,11),
TO_SIGNED(-675,11),
TO_SIGNED(-653,11),
TO_SIGNED(-629,11),
TO_SIGNED(-602,11),
TO_SIGNED(-573,11),
TO_SIGNED(-541,11),
TO_SIGNED(-508,11),
TO_SIGNED(-472,11),
TO_SIGNED(-435,11),
TO_SIGNED(-396,11),
TO_SIGNED(-355,11),
TO_SIGNED(-313,11),
TO_SIGNED(-270,11),
TO_SIGNED(-225,11),
TO_SIGNED(-180,11),
TO_SIGNED(-134,11),
TO_SIGNED(-87,11),
TO_SIGNED(-41,11),
TO_SIGNED(6,11),
TO_SIGNED(53,11),
TO_SIGNED(100,11),
TO_SIGNED(147,11),
TO_SIGNED(192,11),
TO_SIGNED(237,11),
TO_SIGNED(281,11),
TO_SIGNED(324,11),
TO_SIGNED(366,11),
TO_SIGNED(406,11),
TO_SIGNED(445,11),
TO_SIGNED(482,11),
TO_SIGNED(517,11),
TO_SIGNED(550,11),
TO_SIGNED(581,11),
TO_SIGNED(610,11),
TO_SIGNED(636,11),
TO_SIGNED(659,11),
TO_SIGNED(681,11),
TO_SIGNED(699,11),
TO_SIGNED(715,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(712,11),
TO_SIGNED(696,11),
TO_SIGNED(677,11),
TO_SIGNED(656,11),
TO_SIGNED(632,11),
TO_SIGNED(605,11),
TO_SIGNED(576,11),
TO_SIGNED(545,11),
TO_SIGNED(512,11),
TO_SIGNED(476,11),
TO_SIGNED(439,11),
TO_SIGNED(400,11),
TO_SIGNED(360,11),
TO_SIGNED(318,11),
TO_SIGNED(275,11),
TO_SIGNED(230,11),
TO_SIGNED(185,11),
TO_SIGNED(139,11),
TO_SIGNED(93,11),
TO_SIGNED(46,11),
TO_SIGNED(-1,11),
TO_SIGNED(-48,11),
TO_SIGNED(-95,11),
TO_SIGNED(-141,11),
TO_SIGNED(-187,11),
TO_SIGNED(-232,11),
TO_SIGNED(-276,11),
TO_SIGNED(-320,11),
TO_SIGNED(-362,11),
TO_SIGNED(-402,11),
TO_SIGNED(-441,11),
TO_SIGNED(-478,11),
TO_SIGNED(-513,11),
TO_SIGNED(-547,11),
TO_SIGNED(-578,11),
TO_SIGNED(-606,11),
TO_SIGNED(-633,11),
TO_SIGNED(-657,11),
TO_SIGNED(-678,11),
TO_SIGNED(-697,11),
TO_SIGNED(-713,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-714,11),
TO_SIGNED(-698,11),
TO_SIGNED(-680,11),
TO_SIGNED(-658,11),
TO_SIGNED(-635,11),
TO_SIGNED(-608,11),
TO_SIGNED(-580,11),
TO_SIGNED(-549,11),
TO_SIGNED(-516,11),
TO_SIGNED(-480,11),
TO_SIGNED(-443,11),
TO_SIGNED(-405,11),
TO_SIGNED(-364,11),
TO_SIGNED(-323,11),
TO_SIGNED(-279,11),
TO_SIGNED(-235,11),
TO_SIGNED(-190,11),
TO_SIGNED(-144,11),
TO_SIGNED(-98,11),
TO_SIGNED(-51,11),
TO_SIGNED(-4,11),
TO_SIGNED(43,11),
TO_SIGNED(90,11),
TO_SIGNED(136,11),
TO_SIGNED(182,11),
TO_SIGNED(227,11),
TO_SIGNED(272,11),
TO_SIGNED(315,11),
TO_SIGNED(357,11),
TO_SIGNED(397,11),
TO_SIGNED(437,11),
TO_SIGNED(474,11),
TO_SIGNED(509,11),
TO_SIGNED(543,11),
TO_SIGNED(574,11),
TO_SIGNED(603,11),
TO_SIGNED(630,11),
TO_SIGNED(654,11),
TO_SIGNED(676,11),
TO_SIGNED(695,11),
TO_SIGNED(711,11),
TO_SIGNED(725,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(716,11),
TO_SIGNED(700,11),
TO_SIGNED(682,11),
TO_SIGNED(661,11),
TO_SIGNED(637,11),
TO_SIGNED(611,11),
TO_SIGNED(583,11),
TO_SIGNED(552,11),
TO_SIGNED(519,11),
TO_SIGNED(485,11),
TO_SIGNED(448,11),
TO_SIGNED(409,11),
TO_SIGNED(369,11),
TO_SIGNED(327,11),
TO_SIGNED(284,11),
TO_SIGNED(240,11),
TO_SIGNED(195,11),
TO_SIGNED(150,11),
TO_SIGNED(103,11),
TO_SIGNED(57,11),
TO_SIGNED(10,11),
TO_SIGNED(-37,11),
TO_SIGNED(-84,11),
TO_SIGNED(-131,11),
TO_SIGNED(-177,11),
TO_SIGNED(-222,11),
TO_SIGNED(-267,11),
TO_SIGNED(-310,11),
TO_SIGNED(-352,11),
TO_SIGNED(-393,11),
TO_SIGNED(-432,11),
TO_SIGNED(-470,11),
TO_SIGNED(-505,11),
TO_SIGNED(-539,11),
TO_SIGNED(-571,11),
TO_SIGNED(-600,11),
TO_SIGNED(-627,11),
TO_SIGNED(-652,11),
TO_SIGNED(-674,11),
TO_SIGNED(-693,11),
TO_SIGNED(-710,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-702,11),
TO_SIGNED(-684,11),
TO_SIGNED(-663,11),
TO_SIGNED(-640,11),
TO_SIGNED(-615,11),
TO_SIGNED(-586,11),
TO_SIGNED(-556,11),
TO_SIGNED(-523,11),
TO_SIGNED(-489,11),
TO_SIGNED(-452,11),
TO_SIGNED(-414,11),
TO_SIGNED(-374,11),
TO_SIGNED(-332,11),
TO_SIGNED(-289,11),
TO_SIGNED(-245,11),
TO_SIGNED(-201,11),
TO_SIGNED(-155,11),
TO_SIGNED(-109,11),
TO_SIGNED(-62,11),
TO_SIGNED(-15,11),
TO_SIGNED(32,11),
TO_SIGNED(79,11),
TO_SIGNED(125,11),
TO_SIGNED(172,11),
TO_SIGNED(217,11),
TO_SIGNED(262,11),
TO_SIGNED(305,11),
TO_SIGNED(347,11),
TO_SIGNED(388,11),
TO_SIGNED(428,11),
TO_SIGNED(466,11),
TO_SIGNED(501,11),
TO_SIGNED(535,11),
TO_SIGNED(567,11),
TO_SIGNED(597,11),
TO_SIGNED(624,11),
TO_SIGNED(649,11),
TO_SIGNED(671,11),
TO_SIGNED(691,11),
TO_SIGNED(708,11),
TO_SIGNED(722,11),
TO_SIGNED(733,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(704,11),
TO_SIGNED(686,11),
TO_SIGNED(666,11),
TO_SIGNED(643,11),
TO_SIGNED(618,11),
TO_SIGNED(590,11),
TO_SIGNED(559,11),
TO_SIGNED(527,11),
TO_SIGNED(493,11),
TO_SIGNED(456,11),
TO_SIGNED(418,11),
TO_SIGNED(378,11),
TO_SIGNED(337,11),
TO_SIGNED(294,11),
TO_SIGNED(250,11),
TO_SIGNED(206,11),
TO_SIGNED(160,11),
TO_SIGNED(114,11),
TO_SIGNED(67,11),
TO_SIGNED(20,11),
TO_SIGNED(-27,11),
TO_SIGNED(-74,11),
TO_SIGNED(-120,11),
TO_SIGNED(-166,11),
TO_SIGNED(-212,11),
TO_SIGNED(-257,11),
TO_SIGNED(-300,11),
TO_SIGNED(-343,11),
TO_SIGNED(-384,11),
TO_SIGNED(-423,11),
TO_SIGNED(-461,11),
TO_SIGNED(-497,11),
TO_SIGNED(-532,11),
TO_SIGNED(-564,11),
TO_SIGNED(-594,11),
TO_SIGNED(-621,11),
TO_SIGNED(-646,11),
TO_SIGNED(-669,11),
TO_SIGNED(-689,11),
TO_SIGNED(-706,11),
TO_SIGNED(-721,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-720,11),
TO_SIGNED(-706,11),
TO_SIGNED(-688,11),
TO_SIGNED(-668,11),
TO_SIGNED(-646,11),
TO_SIGNED(-621,11),
TO_SIGNED(-593,11),
TO_SIGNED(-563,11),
TO_SIGNED(-531,11),
TO_SIGNED(-497,11),
TO_SIGNED(-460,11),
TO_SIGNED(-422,11),
TO_SIGNED(-383,11),
TO_SIGNED(-342,11),
TO_SIGNED(-299,11),
TO_SIGNED(-256,11),
TO_SIGNED(-211,11),
TO_SIGNED(-165,11),
TO_SIGNED(-119,11),
TO_SIGNED(-73,11),
TO_SIGNED(-26,11),
TO_SIGNED(21,11),
TO_SIGNED(68,11),
TO_SIGNED(115,11),
TO_SIGNED(161,11),
TO_SIGNED(207,11),
TO_SIGNED(251,11),
TO_SIGNED(295,11),
TO_SIGNED(338,11),
TO_SIGNED(379,11),
TO_SIGNED(419,11),
TO_SIGNED(457,11),
TO_SIGNED(493,11),
TO_SIGNED(528,11),
TO_SIGNED(560,11),
TO_SIGNED(590,11),
TO_SIGNED(618,11),
TO_SIGNED(644,11),
TO_SIGNED(666,11),
TO_SIGNED(687,11),
TO_SIGNED(704,11),
TO_SIGNED(719,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(671,11),
TO_SIGNED(648,11),
TO_SIGNED(624,11),
TO_SIGNED(596,11),
TO_SIGNED(567,11),
TO_SIGNED(535,11),
TO_SIGNED(501,11),
TO_SIGNED(465,11),
TO_SIGNED(427,11),
TO_SIGNED(387,11),
TO_SIGNED(346,11),
TO_SIGNED(304,11),
TO_SIGNED(261,11),
TO_SIGNED(216,11),
TO_SIGNED(171,11),
TO_SIGNED(124,11),
TO_SIGNED(78,11),
TO_SIGNED(31,11),
TO_SIGNED(-16,11),
TO_SIGNED(-63,11),
TO_SIGNED(-110,11),
TO_SIGNED(-156,11),
TO_SIGNED(-202,11),
TO_SIGNED(-246,11),
TO_SIGNED(-290,11),
TO_SIGNED(-333,11),
TO_SIGNED(-375,11),
TO_SIGNED(-415,11),
TO_SIGNED(-453,11),
TO_SIGNED(-489,11),
TO_SIGNED(-524,11),
TO_SIGNED(-557,11),
TO_SIGNED(-587,11),
TO_SIGNED(-615,11),
TO_SIGNED(-641,11),
TO_SIGNED(-664,11),
TO_SIGNED(-685,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-730,11),
TO_SIGNED(-739,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-693,11),
TO_SIGNED(-673,11),
TO_SIGNED(-651,11),
TO_SIGNED(-627,11),
TO_SIGNED(-599,11),
TO_SIGNED(-570,11),
TO_SIGNED(-538,11),
TO_SIGNED(-505,11),
TO_SIGNED(-469,11),
TO_SIGNED(-431,11),
TO_SIGNED(-392,11),
TO_SIGNED(-351,11),
TO_SIGNED(-309,11),
TO_SIGNED(-266,11),
TO_SIGNED(-221,11),
TO_SIGNED(-176,11),
TO_SIGNED(-130,11),
TO_SIGNED(-83,11),
TO_SIGNED(-36,11),
TO_SIGNED(11,11),
TO_SIGNED(58,11),
TO_SIGNED(104,11),
TO_SIGNED(151,11),
TO_SIGNED(196,11),
TO_SIGNED(241,11),
TO_SIGNED(285,11),
TO_SIGNED(328,11),
TO_SIGNED(370,11),
TO_SIGNED(410,11),
TO_SIGNED(449,11),
TO_SIGNED(485,11),
TO_SIGNED(520,11),
TO_SIGNED(553,11),
TO_SIGNED(584,11),
TO_SIGNED(612,11),
TO_SIGNED(638,11),
TO_SIGNED(661,11),
TO_SIGNED(682,11),
TO_SIGNED(700,11),
TO_SIGNED(716,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(725,11),
TO_SIGNED(711,11),
TO_SIGNED(695,11),
TO_SIGNED(675,11),
TO_SIGNED(654,11),
TO_SIGNED(629,11),
TO_SIGNED(603,11),
TO_SIGNED(574,11),
TO_SIGNED(542,11),
TO_SIGNED(509,11),
TO_SIGNED(473,11),
TO_SIGNED(436,11),
TO_SIGNED(397,11),
TO_SIGNED(356,11),
TO_SIGNED(314,11),
TO_SIGNED(271,11),
TO_SIGNED(226,11),
TO_SIGNED(181,11),
TO_SIGNED(135,11),
TO_SIGNED(88,11),
TO_SIGNED(42,11),
TO_SIGNED(-5,11),
TO_SIGNED(-52,11),
TO_SIGNED(-99,11),
TO_SIGNED(-145,11),
TO_SIGNED(-191,11),
TO_SIGNED(-236,11),
TO_SIGNED(-280,11),
TO_SIGNED(-323,11),
TO_SIGNED(-365,11),
TO_SIGNED(-406,11),
TO_SIGNED(-444,11),
TO_SIGNED(-481,11),
TO_SIGNED(-516,11),
TO_SIGNED(-549,11),
TO_SIGNED(-580,11),
TO_SIGNED(-609,11),
TO_SIGNED(-635,11),
TO_SIGNED(-659,11),
TO_SIGNED(-680,11),
TO_SIGNED(-699,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-736,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-678,11),
TO_SIGNED(-656,11),
TO_SIGNED(-632,11),
TO_SIGNED(-606,11),
TO_SIGNED(-577,11),
TO_SIGNED(-546,11),
TO_SIGNED(-512,11),
TO_SIGNED(-477,11),
TO_SIGNED(-440,11),
TO_SIGNED(-401,11),
TO_SIGNED(-361,11),
TO_SIGNED(-319,11),
TO_SIGNED(-275,11),
TO_SIGNED(-231,11),
TO_SIGNED(-186,11),
TO_SIGNED(-140,11),
TO_SIGNED(-94,11),
TO_SIGNED(-47,11),
TO_SIGNED(0,11),
TO_SIGNED(47,11),
TO_SIGNED(94,11),
TO_SIGNED(140,11),
TO_SIGNED(186,11),
TO_SIGNED(231,11),
TO_SIGNED(275,11),
TO_SIGNED(319,11),
TO_SIGNED(361,11),
TO_SIGNED(401,11),
TO_SIGNED(440,11),
TO_SIGNED(477,11),
TO_SIGNED(512,11),
TO_SIGNED(546,11),
TO_SIGNED(577,11),
TO_SIGNED(606,11),
TO_SIGNED(632,11),
TO_SIGNED(656,11),
TO_SIGNED(678,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(736,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(699,11),
TO_SIGNED(680,11),
TO_SIGNED(659,11),
TO_SIGNED(635,11),
TO_SIGNED(609,11),
TO_SIGNED(580,11),
TO_SIGNED(549,11),
TO_SIGNED(516,11),
TO_SIGNED(481,11),
TO_SIGNED(444,11),
TO_SIGNED(406,11),
TO_SIGNED(365,11),
TO_SIGNED(323,11),
TO_SIGNED(280,11),
TO_SIGNED(236,11),
TO_SIGNED(191,11),
TO_SIGNED(145,11),
TO_SIGNED(99,11),
TO_SIGNED(52,11),
TO_SIGNED(5,11),
TO_SIGNED(-42,11),
TO_SIGNED(-88,11),
TO_SIGNED(-135,11),
TO_SIGNED(-181,11),
TO_SIGNED(-226,11),
TO_SIGNED(-271,11),
TO_SIGNED(-314,11),
TO_SIGNED(-356,11),
TO_SIGNED(-397,11),
TO_SIGNED(-436,11),
TO_SIGNED(-473,11),
TO_SIGNED(-509,11),
TO_SIGNED(-542,11),
TO_SIGNED(-574,11),
TO_SIGNED(-603,11),
TO_SIGNED(-629,11),
TO_SIGNED(-654,11),
TO_SIGNED(-675,11),
TO_SIGNED(-695,11),
TO_SIGNED(-711,11),
TO_SIGNED(-725,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-716,11),
TO_SIGNED(-700,11),
TO_SIGNED(-682,11),
TO_SIGNED(-661,11),
TO_SIGNED(-638,11),
TO_SIGNED(-612,11),
TO_SIGNED(-584,11),
TO_SIGNED(-553,11),
TO_SIGNED(-520,11),
TO_SIGNED(-485,11),
TO_SIGNED(-449,11),
TO_SIGNED(-410,11),
TO_SIGNED(-370,11),
TO_SIGNED(-328,11),
TO_SIGNED(-285,11),
TO_SIGNED(-241,11),
TO_SIGNED(-196,11),
TO_SIGNED(-151,11),
TO_SIGNED(-104,11),
TO_SIGNED(-58,11),
TO_SIGNED(-11,11),
TO_SIGNED(36,11),
TO_SIGNED(83,11),
TO_SIGNED(130,11),
TO_SIGNED(176,11),
TO_SIGNED(221,11),
TO_SIGNED(266,11),
TO_SIGNED(309,11),
TO_SIGNED(351,11),
TO_SIGNED(392,11),
TO_SIGNED(431,11),
TO_SIGNED(469,11),
TO_SIGNED(505,11),
TO_SIGNED(538,11),
TO_SIGNED(570,11),
TO_SIGNED(599,11),
TO_SIGNED(627,11),
TO_SIGNED(651,11),
TO_SIGNED(673,11),
TO_SIGNED(693,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(739,11),
TO_SIGNED(730,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(685,11),
TO_SIGNED(664,11),
TO_SIGNED(641,11),
TO_SIGNED(615,11),
TO_SIGNED(587,11),
TO_SIGNED(557,11),
TO_SIGNED(524,11),
TO_SIGNED(489,11),
TO_SIGNED(453,11),
TO_SIGNED(415,11),
TO_SIGNED(375,11),
TO_SIGNED(333,11),
TO_SIGNED(290,11),
TO_SIGNED(246,11),
TO_SIGNED(202,11),
TO_SIGNED(156,11),
TO_SIGNED(110,11),
TO_SIGNED(63,11),
TO_SIGNED(16,11),
TO_SIGNED(-31,11),
TO_SIGNED(-78,11),
TO_SIGNED(-124,11),
TO_SIGNED(-171,11),
TO_SIGNED(-216,11),
TO_SIGNED(-261,11),
TO_SIGNED(-304,11),
TO_SIGNED(-346,11),
TO_SIGNED(-387,11),
TO_SIGNED(-427,11),
TO_SIGNED(-465,11),
TO_SIGNED(-501,11),
TO_SIGNED(-535,11),
TO_SIGNED(-567,11),
TO_SIGNED(-596,11),
TO_SIGNED(-624,11),
TO_SIGNED(-648,11),
TO_SIGNED(-671,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-719,11),
TO_SIGNED(-704,11),
TO_SIGNED(-687,11),
TO_SIGNED(-666,11),
TO_SIGNED(-644,11),
TO_SIGNED(-618,11),
TO_SIGNED(-590,11),
TO_SIGNED(-560,11),
TO_SIGNED(-528,11),
TO_SIGNED(-493,11),
TO_SIGNED(-457,11),
TO_SIGNED(-419,11),
TO_SIGNED(-379,11),
TO_SIGNED(-338,11),
TO_SIGNED(-295,11),
TO_SIGNED(-251,11),
TO_SIGNED(-207,11),
TO_SIGNED(-161,11),
TO_SIGNED(-115,11),
TO_SIGNED(-68,11),
TO_SIGNED(-21,11),
TO_SIGNED(26,11),
TO_SIGNED(73,11),
TO_SIGNED(119,11),
TO_SIGNED(165,11),
TO_SIGNED(211,11),
TO_SIGNED(256,11),
TO_SIGNED(299,11),
TO_SIGNED(342,11),
TO_SIGNED(383,11),
TO_SIGNED(422,11),
TO_SIGNED(460,11),
TO_SIGNED(497,11),
TO_SIGNED(531,11),
TO_SIGNED(563,11),
TO_SIGNED(593,11),
TO_SIGNED(621,11),
TO_SIGNED(646,11),
TO_SIGNED(668,11),
TO_SIGNED(688,11),
TO_SIGNED(706,11),
TO_SIGNED(720,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(721,11),
TO_SIGNED(706,11),
TO_SIGNED(689,11),
TO_SIGNED(669,11),
TO_SIGNED(646,11),
TO_SIGNED(621,11),
TO_SIGNED(594,11),
TO_SIGNED(564,11),
TO_SIGNED(532,11),
TO_SIGNED(497,11),
TO_SIGNED(461,11),
TO_SIGNED(423,11),
TO_SIGNED(384,11),
TO_SIGNED(343,11),
TO_SIGNED(300,11),
TO_SIGNED(257,11),
TO_SIGNED(212,11),
TO_SIGNED(166,11),
TO_SIGNED(120,11),
TO_SIGNED(74,11),
TO_SIGNED(27,11),
TO_SIGNED(-20,11),
TO_SIGNED(-67,11),
TO_SIGNED(-114,11),
TO_SIGNED(-160,11),
TO_SIGNED(-206,11),
TO_SIGNED(-250,11),
TO_SIGNED(-294,11),
TO_SIGNED(-337,11),
TO_SIGNED(-378,11),
TO_SIGNED(-418,11),
TO_SIGNED(-456,11),
TO_SIGNED(-493,11),
TO_SIGNED(-527,11),
TO_SIGNED(-559,11),
TO_SIGNED(-590,11),
TO_SIGNED(-618,11),
TO_SIGNED(-643,11),
TO_SIGNED(-666,11),
TO_SIGNED(-686,11),
TO_SIGNED(-704,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-733,11),
TO_SIGNED(-722,11),
TO_SIGNED(-708,11),
TO_SIGNED(-691,11),
TO_SIGNED(-671,11),
TO_SIGNED(-649,11),
TO_SIGNED(-624,11),
TO_SIGNED(-597,11),
TO_SIGNED(-567,11),
TO_SIGNED(-535,11),
TO_SIGNED(-501,11),
TO_SIGNED(-466,11),
TO_SIGNED(-428,11),
TO_SIGNED(-388,11),
TO_SIGNED(-347,11),
TO_SIGNED(-305,11),
TO_SIGNED(-262,11),
TO_SIGNED(-217,11),
TO_SIGNED(-172,11),
TO_SIGNED(-125,11),
TO_SIGNED(-79,11),
TO_SIGNED(-32,11),
TO_SIGNED(15,11),
TO_SIGNED(62,11),
TO_SIGNED(109,11),
TO_SIGNED(155,11),
TO_SIGNED(201,11),
TO_SIGNED(245,11),
TO_SIGNED(289,11),
TO_SIGNED(332,11),
TO_SIGNED(374,11),
TO_SIGNED(414,11),
TO_SIGNED(452,11),
TO_SIGNED(489,11),
TO_SIGNED(523,11),
TO_SIGNED(556,11),
TO_SIGNED(586,11),
TO_SIGNED(615,11),
TO_SIGNED(640,11),
TO_SIGNED(663,11),
TO_SIGNED(684,11),
TO_SIGNED(702,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(710,11),
TO_SIGNED(693,11),
TO_SIGNED(674,11),
TO_SIGNED(652,11),
TO_SIGNED(627,11),
TO_SIGNED(600,11),
TO_SIGNED(571,11),
TO_SIGNED(539,11),
TO_SIGNED(505,11),
TO_SIGNED(470,11),
TO_SIGNED(432,11),
TO_SIGNED(393,11),
TO_SIGNED(352,11),
TO_SIGNED(310,11),
TO_SIGNED(267,11),
TO_SIGNED(222,11),
TO_SIGNED(177,11),
TO_SIGNED(131,11),
TO_SIGNED(84,11),
TO_SIGNED(37,11),
TO_SIGNED(-10,11),
TO_SIGNED(-57,11),
TO_SIGNED(-103,11),
TO_SIGNED(-150,11),
TO_SIGNED(-195,11),
TO_SIGNED(-240,11),
TO_SIGNED(-284,11),
TO_SIGNED(-327,11),
TO_SIGNED(-369,11),
TO_SIGNED(-409,11),
TO_SIGNED(-448,11),
TO_SIGNED(-485,11),
TO_SIGNED(-519,11),
TO_SIGNED(-552,11),
TO_SIGNED(-583,11),
TO_SIGNED(-611,11),
TO_SIGNED(-637,11),
TO_SIGNED(-661,11),
TO_SIGNED(-682,11),
TO_SIGNED(-700,11),
TO_SIGNED(-716,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-725,11),
TO_SIGNED(-711,11),
TO_SIGNED(-695,11),
TO_SIGNED(-676,11),
TO_SIGNED(-654,11),
TO_SIGNED(-630,11),
TO_SIGNED(-603,11),
TO_SIGNED(-574,11),
TO_SIGNED(-543,11),
TO_SIGNED(-509,11),
TO_SIGNED(-474,11),
TO_SIGNED(-437,11),
TO_SIGNED(-397,11),
TO_SIGNED(-357,11),
TO_SIGNED(-315,11),
TO_SIGNED(-272,11),
TO_SIGNED(-227,11),
TO_SIGNED(-182,11),
TO_SIGNED(-136,11),
TO_SIGNED(-90,11),
TO_SIGNED(-43,11),
TO_SIGNED(4,11),
TO_SIGNED(51,11),
TO_SIGNED(98,11),
TO_SIGNED(144,11),
TO_SIGNED(190,11),
TO_SIGNED(235,11),
TO_SIGNED(279,11),
TO_SIGNED(323,11),
TO_SIGNED(364,11),
TO_SIGNED(405,11),
TO_SIGNED(443,11),
TO_SIGNED(480,11),
TO_SIGNED(516,11),
TO_SIGNED(549,11),
TO_SIGNED(580,11),
TO_SIGNED(608,11),
TO_SIGNED(635,11),
TO_SIGNED(658,11),
TO_SIGNED(680,11),
TO_SIGNED(698,11),
TO_SIGNED(714,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(713,11),
TO_SIGNED(697,11),
TO_SIGNED(678,11),
TO_SIGNED(657,11),
TO_SIGNED(633,11),
TO_SIGNED(606,11),
TO_SIGNED(578,11),
TO_SIGNED(547,11),
TO_SIGNED(513,11),
TO_SIGNED(478,11),
TO_SIGNED(441,11),
TO_SIGNED(402,11),
TO_SIGNED(362,11),
TO_SIGNED(320,11),
TO_SIGNED(276,11),
TO_SIGNED(232,11),
TO_SIGNED(187,11),
TO_SIGNED(141,11),
TO_SIGNED(95,11),
TO_SIGNED(48,11),
TO_SIGNED(1,11),
TO_SIGNED(-46,11),
TO_SIGNED(-93,11),
TO_SIGNED(-139,11),
TO_SIGNED(-185,11),
TO_SIGNED(-230,11),
TO_SIGNED(-275,11),
TO_SIGNED(-318,11),
TO_SIGNED(-360,11),
TO_SIGNED(-400,11),
TO_SIGNED(-439,11),
TO_SIGNED(-476,11),
TO_SIGNED(-512,11),
TO_SIGNED(-545,11),
TO_SIGNED(-576,11),
TO_SIGNED(-605,11),
TO_SIGNED(-632,11),
TO_SIGNED(-656,11),
TO_SIGNED(-677,11),
TO_SIGNED(-696,11),
TO_SIGNED(-712,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-715,11),
TO_SIGNED(-699,11),
TO_SIGNED(-681,11),
TO_SIGNED(-659,11),
TO_SIGNED(-636,11),
TO_SIGNED(-610,11),
TO_SIGNED(-581,11),
TO_SIGNED(-550,11),
TO_SIGNED(-517,11),
TO_SIGNED(-482,11),
TO_SIGNED(-445,11),
TO_SIGNED(-406,11),
TO_SIGNED(-366,11),
TO_SIGNED(-324,11),
TO_SIGNED(-281,11),
TO_SIGNED(-237,11),
TO_SIGNED(-192,11),
TO_SIGNED(-147,11),
TO_SIGNED(-100,11),
TO_SIGNED(-53,11),
TO_SIGNED(-6,11),
TO_SIGNED(41,11),
TO_SIGNED(87,11),
TO_SIGNED(134,11),
TO_SIGNED(180,11),
TO_SIGNED(225,11),
TO_SIGNED(270,11),
TO_SIGNED(313,11),
TO_SIGNED(355,11),
TO_SIGNED(396,11),
TO_SIGNED(435,11),
TO_SIGNED(472,11),
TO_SIGNED(508,11),
TO_SIGNED(541,11),
TO_SIGNED(573,11),
TO_SIGNED(602,11),
TO_SIGNED(629,11),
TO_SIGNED(653,11),
TO_SIGNED(675,11),
TO_SIGNED(694,11),
TO_SIGNED(711,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(729,11),
TO_SIGNED(716,11),
TO_SIGNED(701,11),
TO_SIGNED(683,11),
TO_SIGNED(662,11),
TO_SIGNED(639,11),
TO_SIGNED(613,11),
TO_SIGNED(584,11),
TO_SIGNED(554,11),
TO_SIGNED(521,11),
TO_SIGNED(486,11),
TO_SIGNED(449,11),
TO_SIGNED(411,11),
TO_SIGNED(371,11),
TO_SIGNED(329,11),
TO_SIGNED(286,11),
TO_SIGNED(242,11),
TO_SIGNED(197,11),
TO_SIGNED(152,11),
TO_SIGNED(105,11),
TO_SIGNED(59,11),
TO_SIGNED(12,11),
TO_SIGNED(-35,11),
TO_SIGNED(-82,11),
TO_SIGNED(-129,11),
TO_SIGNED(-175,11),
TO_SIGNED(-220,11),
TO_SIGNED(-265,11),
TO_SIGNED(-308,11),
TO_SIGNED(-350,11),
TO_SIGNED(-391,11),
TO_SIGNED(-430,11),
TO_SIGNED(-468,11),
TO_SIGNED(-504,11),
TO_SIGNED(-538,11),
TO_SIGNED(-569,11),
TO_SIGNED(-599,11),
TO_SIGNED(-626,11),
TO_SIGNED(-651,11),
TO_SIGNED(-673,11),
TO_SIGNED(-692,11),
TO_SIGNED(-709,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-685,11),
TO_SIGNED(-664,11),
TO_SIGNED(-641,11),
TO_SIGNED(-616,11),
TO_SIGNED(-588,11),
TO_SIGNED(-557,11),
TO_SIGNED(-525,11),
TO_SIGNED(-490,11),
TO_SIGNED(-454,11),
TO_SIGNED(-415,11),
TO_SIGNED(-375,11),
TO_SIGNED(-334,11),
TO_SIGNED(-291,11),
TO_SIGNED(-247,11),
TO_SIGNED(-203,11),
TO_SIGNED(-157,11),
TO_SIGNED(-111,11),
TO_SIGNED(-64,11),
TO_SIGNED(-17,11),
TO_SIGNED(30,11),
TO_SIGNED(77,11),
TO_SIGNED(123,11),
TO_SIGNED(169,11),
TO_SIGNED(215,11),
TO_SIGNED(260,11),
TO_SIGNED(303,11),
TO_SIGNED(345,11),
TO_SIGNED(387,11),
TO_SIGNED(426,11),
TO_SIGNED(464,11),
TO_SIGNED(500,11),
TO_SIGNED(534,11),
TO_SIGNED(566,11),
TO_SIGNED(596,11),
TO_SIGNED(623,11),
TO_SIGNED(648,11),
TO_SIGNED(670,11),
TO_SIGNED(690,11),
TO_SIGNED(707,11),
TO_SIGNED(721,11),
TO_SIGNED(733,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(705,11),
TO_SIGNED(687,11),
TO_SIGNED(667,11),
TO_SIGNED(644,11),
TO_SIGNED(619,11),
TO_SIGNED(591,11),
TO_SIGNED(561,11),
TO_SIGNED(529,11),
TO_SIGNED(494,11),
TO_SIGNED(458,11),
TO_SIGNED(420,11),
TO_SIGNED(380,11),
TO_SIGNED(339,11),
TO_SIGNED(296,11),
TO_SIGNED(252,11),
TO_SIGNED(208,11),
TO_SIGNED(162,11),
TO_SIGNED(116,11),
TO_SIGNED(69,11),
TO_SIGNED(22,11),
TO_SIGNED(-25,11),
TO_SIGNED(-71,11),
TO_SIGNED(-118,11),
TO_SIGNED(-164,11),
TO_SIGNED(-210,11),
TO_SIGNED(-255,11),
TO_SIGNED(-298,11),
TO_SIGNED(-341,11),
TO_SIGNED(-382,11),
TO_SIGNED(-422,11),
TO_SIGNED(-460,11),
TO_SIGNED(-496,11),
TO_SIGNED(-530,11),
TO_SIGNED(-562,11),
TO_SIGNED(-592,11),
TO_SIGNED(-620,11),
TO_SIGNED(-645,11),
TO_SIGNED(-668,11),
TO_SIGNED(-688,11),
TO_SIGNED(-705,11),
TO_SIGNED(-720,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-721,11),
TO_SIGNED(-706,11),
TO_SIGNED(-689,11),
TO_SIGNED(-669,11),
TO_SIGNED(-647,11),
TO_SIGNED(-622,11),
TO_SIGNED(-594,11),
TO_SIGNED(-564,11),
TO_SIGNED(-532,11),
TO_SIGNED(-498,11),
TO_SIGNED(-462,11),
TO_SIGNED(-424,11),
TO_SIGNED(-385,11),
TO_SIGNED(-344,11),
TO_SIGNED(-301,11),
TO_SIGNED(-258,11),
TO_SIGNED(-213,11),
TO_SIGNED(-167,11),
TO_SIGNED(-121,11),
TO_SIGNED(-75,11),
TO_SIGNED(-28,11),
TO_SIGNED(19,11),
TO_SIGNED(66,11),
TO_SIGNED(113,11),
TO_SIGNED(159,11),
TO_SIGNED(205,11),
TO_SIGNED(249,11),
TO_SIGNED(293,11),
TO_SIGNED(336,11),
TO_SIGNED(377,11),
TO_SIGNED(417,11),
TO_SIGNED(455,11),
TO_SIGNED(492,11),
TO_SIGNED(526,11),
TO_SIGNED(559,11),
TO_SIGNED(589,11),
TO_SIGNED(617,11),
TO_SIGNED(642,11),
TO_SIGNED(665,11),
TO_SIGNED(686,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(708,11),
TO_SIGNED(691,11),
TO_SIGNED(672,11),
TO_SIGNED(650,11),
TO_SIGNED(625,11),
TO_SIGNED(598,11),
TO_SIGNED(568,11),
TO_SIGNED(536,11),
TO_SIGNED(502,11),
TO_SIGNED(466,11),
TO_SIGNED(429,11),
TO_SIGNED(389,11),
TO_SIGNED(348,11),
TO_SIGNED(306,11),
TO_SIGNED(263,11),
TO_SIGNED(218,11),
TO_SIGNED(173,11),
TO_SIGNED(127,11),
TO_SIGNED(80,11),
TO_SIGNED(33,11),
TO_SIGNED(-14,11),
TO_SIGNED(-61,11),
TO_SIGNED(-108,11),
TO_SIGNED(-154,11),
TO_SIGNED(-200,11),
TO_SIGNED(-244,11),
TO_SIGNED(-288,11),
TO_SIGNED(-331,11),
TO_SIGNED(-373,11),
TO_SIGNED(-413,11),
TO_SIGNED(-451,11),
TO_SIGNED(-488,11),
TO_SIGNED(-523,11),
TO_SIGNED(-555,11),
TO_SIGNED(-586,11),
TO_SIGNED(-614,11),
TO_SIGNED(-640,11),
TO_SIGNED(-663,11),
TO_SIGNED(-684,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-729,11),
TO_SIGNED(-739,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-710,11),
TO_SIGNED(-693,11),
TO_SIGNED(-674,11),
TO_SIGNED(-652,11),
TO_SIGNED(-628,11),
TO_SIGNED(-601,11),
TO_SIGNED(-571,11),
TO_SIGNED(-540,11),
TO_SIGNED(-506,11),
TO_SIGNED(-471,11),
TO_SIGNED(-433,11),
TO_SIGNED(-394,11),
TO_SIGNED(-353,11),
TO_SIGNED(-311,11),
TO_SIGNED(-268,11),
TO_SIGNED(-223,11),
TO_SIGNED(-178,11),
TO_SIGNED(-132,11),
TO_SIGNED(-85,11),
TO_SIGNED(-38,11),
TO_SIGNED(9,11),
TO_SIGNED(56,11),
TO_SIGNED(102,11),
TO_SIGNED(149,11),
TO_SIGNED(194,11),
TO_SIGNED(239,11),
TO_SIGNED(283,11),
TO_SIGNED(326,11),
TO_SIGNED(368,11),
TO_SIGNED(408,11),
TO_SIGNED(447,11),
TO_SIGNED(484,11),
TO_SIGNED(519,11),
TO_SIGNED(552,11),
TO_SIGNED(582,11),
TO_SIGNED(611,11),
TO_SIGNED(637,11),
TO_SIGNED(660,11),
TO_SIGNED(681,11),
TO_SIGNED(700,11),
TO_SIGNED(715,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(736,11),
TO_SIGNED(725,11),
TO_SIGNED(712,11),
TO_SIGNED(695,11),
TO_SIGNED(676,11),
TO_SIGNED(655,11),
TO_SIGNED(631,11),
TO_SIGNED(604,11),
TO_SIGNED(575,11),
TO_SIGNED(544,11),
TO_SIGNED(510,11),
TO_SIGNED(475,11),
TO_SIGNED(437,11),
TO_SIGNED(398,11),
TO_SIGNED(358,11),
TO_SIGNED(316,11),
TO_SIGNED(273,11),
TO_SIGNED(228,11),
TO_SIGNED(183,11),
TO_SIGNED(137,11),
TO_SIGNED(91,11),
TO_SIGNED(44,11),
TO_SIGNED(-3,11),
TO_SIGNED(-50,11),
TO_SIGNED(-97,11),
TO_SIGNED(-143,11),
TO_SIGNED(-189,11),
TO_SIGNED(-234,11),
TO_SIGNED(-278,11),
TO_SIGNED(-322,11),
TO_SIGNED(-363,11),
TO_SIGNED(-404,11),
TO_SIGNED(-443,11),
TO_SIGNED(-480,11),
TO_SIGNED(-515,11),
TO_SIGNED(-548,11),
TO_SIGNED(-579,11),
TO_SIGNED(-608,11),
TO_SIGNED(-634,11),
TO_SIGNED(-658,11),
TO_SIGNED(-679,11),
TO_SIGNED(-698,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-679,11),
TO_SIGNED(-657,11),
TO_SIGNED(-633,11),
TO_SIGNED(-607,11),
TO_SIGNED(-578,11),
TO_SIGNED(-547,11),
TO_SIGNED(-514,11),
TO_SIGNED(-479,11),
TO_SIGNED(-442,11),
TO_SIGNED(-403,11),
TO_SIGNED(-362,11),
TO_SIGNED(-321,11),
TO_SIGNED(-277,11),
TO_SIGNED(-233,11),
TO_SIGNED(-188,11),
TO_SIGNED(-142,11),
TO_SIGNED(-96,11),
TO_SIGNED(-49,11),
TO_SIGNED(-2,11),
TO_SIGNED(45,11),
TO_SIGNED(92,11),
TO_SIGNED(138,11),
TO_SIGNED(184,11),
TO_SIGNED(229,11),
TO_SIGNED(274,11),
TO_SIGNED(317,11),
TO_SIGNED(359,11),
TO_SIGNED(399,11),
TO_SIGNED(438,11),
TO_SIGNED(476,11),
TO_SIGNED(511,11),
TO_SIGNED(544,11),
TO_SIGNED(576,11),
TO_SIGNED(605,11),
TO_SIGNED(631,11),
TO_SIGNED(655,11),
TO_SIGNED(677,11),
TO_SIGNED(696,11),
TO_SIGNED(712,11),
TO_SIGNED(725,11),
TO_SIGNED(736,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(715,11),
TO_SIGNED(699,11),
TO_SIGNED(681,11),
TO_SIGNED(660,11),
TO_SIGNED(636,11),
TO_SIGNED(610,11),
TO_SIGNED(582,11),
TO_SIGNED(551,11),
TO_SIGNED(518,11),
TO_SIGNED(483,11),
TO_SIGNED(446,11),
TO_SIGNED(407,11),
TO_SIGNED(367,11),
TO_SIGNED(325,11),
TO_SIGNED(282,11),
TO_SIGNED(238,11),
TO_SIGNED(193,11),
TO_SIGNED(148,11),
TO_SIGNED(101,11),
TO_SIGNED(54,11),
TO_SIGNED(7,11),
TO_SIGNED(-40,11),
TO_SIGNED(-86,11),
TO_SIGNED(-133,11),
TO_SIGNED(-179,11),
TO_SIGNED(-224,11),
TO_SIGNED(-269,11),
TO_SIGNED(-312,11),
TO_SIGNED(-354,11),
TO_SIGNED(-395,11),
TO_SIGNED(-434,11),
TO_SIGNED(-471,11),
TO_SIGNED(-507,11),
TO_SIGNED(-541,11),
TO_SIGNED(-572,11),
TO_SIGNED(-601,11),
TO_SIGNED(-628,11),
TO_SIGNED(-653,11),
TO_SIGNED(-675,11),
TO_SIGNED(-694,11),
TO_SIGNED(-710,11),
TO_SIGNED(-724,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-701,11),
TO_SIGNED(-683,11),
TO_SIGNED(-662,11),
TO_SIGNED(-639,11),
TO_SIGNED(-613,11),
TO_SIGNED(-585,11),
TO_SIGNED(-554,11),
TO_SIGNED(-522,11),
TO_SIGNED(-487,11),
TO_SIGNED(-450,11),
TO_SIGNED(-412,11),
TO_SIGNED(-372,11),
TO_SIGNED(-330,11),
TO_SIGNED(-287,11),
TO_SIGNED(-243,11),
TO_SIGNED(-198,11),
TO_SIGNED(-153,11),
TO_SIGNED(-106,11),
TO_SIGNED(-60,11),
TO_SIGNED(-13,11),
TO_SIGNED(34,11),
TO_SIGNED(81,11),
TO_SIGNED(128,11),
TO_SIGNED(174,11),
TO_SIGNED(219,11),
TO_SIGNED(264,11),
TO_SIGNED(307,11),
TO_SIGNED(349,11),
TO_SIGNED(390,11),
TO_SIGNED(430,11),
TO_SIGNED(467,11),
TO_SIGNED(503,11),
TO_SIGNED(537,11),
TO_SIGNED(569,11),
TO_SIGNED(598,11),
TO_SIGNED(625,11),
TO_SIGNED(650,11),
TO_SIGNED(672,11),
TO_SIGNED(692,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(730,11),
TO_SIGNED(718,11),
TO_SIGNED(703,11),
TO_SIGNED(685,11),
TO_SIGNED(665,11),
TO_SIGNED(642,11),
TO_SIGNED(616,11),
TO_SIGNED(588,11),
TO_SIGNED(558,11),
TO_SIGNED(526,11),
TO_SIGNED(491,11),
TO_SIGNED(455,11),
TO_SIGNED(416,11),
TO_SIGNED(376,11),
TO_SIGNED(335,11),
TO_SIGNED(292,11),
TO_SIGNED(248,11),
TO_SIGNED(204,11),
TO_SIGNED(158,11),
TO_SIGNED(112,11),
TO_SIGNED(65,11),
TO_SIGNED(18,11),
TO_SIGNED(-29,11),
TO_SIGNED(-76,11),
TO_SIGNED(-122,11),
TO_SIGNED(-168,11),
TO_SIGNED(-214,11),
TO_SIGNED(-259,11),
TO_SIGNED(-302,11),
TO_SIGNED(-345,11),
TO_SIGNED(-386,11),
TO_SIGNED(-425,11),
TO_SIGNED(-463,11),
TO_SIGNED(-499,11),
TO_SIGNED(-533,11),
TO_SIGNED(-565,11),
TO_SIGNED(-595,11),
TO_SIGNED(-622,11),
TO_SIGNED(-647,11),
TO_SIGNED(-670,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-721,11),
TO_SIGNED(-733,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-720,11),
TO_SIGNED(-705,11),
TO_SIGNED(-688,11),
TO_SIGNED(-667,11),
TO_SIGNED(-645,11),
TO_SIGNED(-619,11),
TO_SIGNED(-592,11),
TO_SIGNED(-562,11),
TO_SIGNED(-529,11),
TO_SIGNED(-495,11),
TO_SIGNED(-459,11),
TO_SIGNED(-421,11),
TO_SIGNED(-381,11),
TO_SIGNED(-340,11),
TO_SIGNED(-297,11),
TO_SIGNED(-254,11),
TO_SIGNED(-209,11),
TO_SIGNED(-163,11),
TO_SIGNED(-117,11),
TO_SIGNED(-70,11),
TO_SIGNED(-24,11),
TO_SIGNED(24,11),
TO_SIGNED(70,11),
TO_SIGNED(117,11),
TO_SIGNED(163,11),
TO_SIGNED(209,11),
TO_SIGNED(254,11),
TO_SIGNED(297,11),
TO_SIGNED(340,11),
TO_SIGNED(381,11),
TO_SIGNED(421,11),
TO_SIGNED(459,11),
TO_SIGNED(495,11),
TO_SIGNED(529,11),
TO_SIGNED(562,11),
TO_SIGNED(592,11),
TO_SIGNED(619,11),
TO_SIGNED(645,11),
TO_SIGNED(667,11),
TO_SIGNED(688,11),
TO_SIGNED(705,11),
TO_SIGNED(720,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(733,11),
TO_SIGNED(721,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(670,11),
TO_SIGNED(647,11),
TO_SIGNED(622,11),
TO_SIGNED(595,11),
TO_SIGNED(565,11),
TO_SIGNED(533,11),
TO_SIGNED(499,11),
TO_SIGNED(463,11),
TO_SIGNED(425,11),
TO_SIGNED(386,11),
TO_SIGNED(345,11),
TO_SIGNED(302,11),
TO_SIGNED(259,11),
TO_SIGNED(214,11),
TO_SIGNED(168,11),
TO_SIGNED(122,11),
TO_SIGNED(76,11),
TO_SIGNED(29,11),
TO_SIGNED(-18,11),
TO_SIGNED(-65,11),
TO_SIGNED(-112,11),
TO_SIGNED(-158,11),
TO_SIGNED(-204,11),
TO_SIGNED(-248,11),
TO_SIGNED(-292,11),
TO_SIGNED(-335,11),
TO_SIGNED(-376,11),
TO_SIGNED(-416,11),
TO_SIGNED(-455,11),
TO_SIGNED(-491,11),
TO_SIGNED(-526,11),
TO_SIGNED(-558,11),
TO_SIGNED(-588,11),
TO_SIGNED(-616,11),
TO_SIGNED(-642,11),
TO_SIGNED(-665,11),
TO_SIGNED(-685,11),
TO_SIGNED(-703,11),
TO_SIGNED(-718,11),
TO_SIGNED(-730,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-692,11),
TO_SIGNED(-672,11),
TO_SIGNED(-650,11),
TO_SIGNED(-625,11),
TO_SIGNED(-598,11),
TO_SIGNED(-569,11),
TO_SIGNED(-537,11),
TO_SIGNED(-503,11),
TO_SIGNED(-467,11),
TO_SIGNED(-430,11),
TO_SIGNED(-390,11),
TO_SIGNED(-349,11),
TO_SIGNED(-307,11),
TO_SIGNED(-264,11),
TO_SIGNED(-219,11),
TO_SIGNED(-174,11),
TO_SIGNED(-128,11),
TO_SIGNED(-81,11),
TO_SIGNED(-34,11),
TO_SIGNED(13,11),
TO_SIGNED(60,11),
TO_SIGNED(106,11),
TO_SIGNED(153,11),
TO_SIGNED(198,11),
TO_SIGNED(243,11),
TO_SIGNED(287,11),
TO_SIGNED(330,11),
TO_SIGNED(372,11),
TO_SIGNED(412,11),
TO_SIGNED(450,11),
TO_SIGNED(487,11),
TO_SIGNED(522,11),
TO_SIGNED(554,11),
TO_SIGNED(585,11),
TO_SIGNED(613,11),
TO_SIGNED(639,11),
TO_SIGNED(662,11),
TO_SIGNED(683,11),
TO_SIGNED(701,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(724,11),
TO_SIGNED(710,11),
TO_SIGNED(694,11),
TO_SIGNED(675,11),
TO_SIGNED(653,11),
TO_SIGNED(628,11),
TO_SIGNED(601,11),
TO_SIGNED(572,11),
TO_SIGNED(541,11),
TO_SIGNED(507,11),
TO_SIGNED(471,11),
TO_SIGNED(434,11),
TO_SIGNED(395,11),
TO_SIGNED(354,11),
TO_SIGNED(312,11),
TO_SIGNED(269,11),
TO_SIGNED(224,11),
TO_SIGNED(179,11),
TO_SIGNED(133,11),
TO_SIGNED(86,11),
TO_SIGNED(40,11),
TO_SIGNED(-7,11),
TO_SIGNED(-54,11),
TO_SIGNED(-101,11),
TO_SIGNED(-148,11),
TO_SIGNED(-193,11),
TO_SIGNED(-238,11),
TO_SIGNED(-282,11),
TO_SIGNED(-325,11),
TO_SIGNED(-367,11),
TO_SIGNED(-407,11),
TO_SIGNED(-446,11),
TO_SIGNED(-483,11),
TO_SIGNED(-518,11),
TO_SIGNED(-551,11),
TO_SIGNED(-582,11),
TO_SIGNED(-610,11),
TO_SIGNED(-636,11),
TO_SIGNED(-660,11),
TO_SIGNED(-681,11),
TO_SIGNED(-699,11),
TO_SIGNED(-715,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-736,11),
TO_SIGNED(-725,11),
TO_SIGNED(-712,11),
TO_SIGNED(-696,11),
TO_SIGNED(-677,11),
TO_SIGNED(-655,11),
TO_SIGNED(-631,11),
TO_SIGNED(-605,11),
TO_SIGNED(-576,11),
TO_SIGNED(-544,11),
TO_SIGNED(-511,11),
TO_SIGNED(-476,11),
TO_SIGNED(-438,11),
TO_SIGNED(-399,11),
TO_SIGNED(-359,11),
TO_SIGNED(-317,11),
TO_SIGNED(-274,11),
TO_SIGNED(-229,11),
TO_SIGNED(-184,11),
TO_SIGNED(-138,11),
TO_SIGNED(-92,11),
TO_SIGNED(-45,11),
TO_SIGNED(2,11),
TO_SIGNED(49,11),
TO_SIGNED(96,11),
TO_SIGNED(142,11),
TO_SIGNED(188,11),
TO_SIGNED(233,11),
TO_SIGNED(277,11),
TO_SIGNED(321,11),
TO_SIGNED(362,11),
TO_SIGNED(403,11),
TO_SIGNED(442,11),
TO_SIGNED(479,11),
TO_SIGNED(514,11),
TO_SIGNED(547,11),
TO_SIGNED(578,11),
TO_SIGNED(607,11),
TO_SIGNED(633,11),
TO_SIGNED(657,11),
TO_SIGNED(679,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(698,11),
TO_SIGNED(679,11),
TO_SIGNED(658,11),
TO_SIGNED(634,11),
TO_SIGNED(608,11),
TO_SIGNED(579,11),
TO_SIGNED(548,11),
TO_SIGNED(515,11),
TO_SIGNED(480,11),
TO_SIGNED(443,11),
TO_SIGNED(404,11),
TO_SIGNED(363,11),
TO_SIGNED(322,11),
TO_SIGNED(278,11),
TO_SIGNED(234,11),
TO_SIGNED(189,11),
TO_SIGNED(143,11),
TO_SIGNED(97,11),
TO_SIGNED(50,11),
TO_SIGNED(3,11),
TO_SIGNED(-44,11),
TO_SIGNED(-91,11),
TO_SIGNED(-137,11),
TO_SIGNED(-183,11),
TO_SIGNED(-228,11),
TO_SIGNED(-273,11),
TO_SIGNED(-316,11),
TO_SIGNED(-358,11),
TO_SIGNED(-398,11),
TO_SIGNED(-437,11),
TO_SIGNED(-475,11),
TO_SIGNED(-510,11),
TO_SIGNED(-544,11),
TO_SIGNED(-575,11),
TO_SIGNED(-604,11),
TO_SIGNED(-631,11),
TO_SIGNED(-655,11),
TO_SIGNED(-676,11),
TO_SIGNED(-695,11),
TO_SIGNED(-712,11),
TO_SIGNED(-725,11),
TO_SIGNED(-736,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-715,11),
TO_SIGNED(-700,11),
TO_SIGNED(-681,11),
TO_SIGNED(-660,11),
TO_SIGNED(-637,11),
TO_SIGNED(-611,11),
TO_SIGNED(-582,11),
TO_SIGNED(-552,11),
TO_SIGNED(-519,11),
TO_SIGNED(-484,11),
TO_SIGNED(-447,11),
TO_SIGNED(-408,11),
TO_SIGNED(-368,11),
TO_SIGNED(-326,11),
TO_SIGNED(-283,11),
TO_SIGNED(-239,11),
TO_SIGNED(-194,11),
TO_SIGNED(-149,11),
TO_SIGNED(-102,11),
TO_SIGNED(-56,11),
TO_SIGNED(-9,11),
TO_SIGNED(38,11),
TO_SIGNED(85,11),
TO_SIGNED(132,11),
TO_SIGNED(178,11),
TO_SIGNED(223,11),
TO_SIGNED(268,11),
TO_SIGNED(311,11),
TO_SIGNED(353,11),
TO_SIGNED(394,11),
TO_SIGNED(433,11),
TO_SIGNED(471,11),
TO_SIGNED(506,11),
TO_SIGNED(540,11),
TO_SIGNED(571,11),
TO_SIGNED(601,11),
TO_SIGNED(628,11),
TO_SIGNED(652,11),
TO_SIGNED(674,11),
TO_SIGNED(693,11),
TO_SIGNED(710,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(739,11),
TO_SIGNED(729,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(684,11),
TO_SIGNED(663,11),
TO_SIGNED(640,11),
TO_SIGNED(614,11),
TO_SIGNED(586,11),
TO_SIGNED(555,11),
TO_SIGNED(523,11),
TO_SIGNED(488,11),
TO_SIGNED(451,11),
TO_SIGNED(413,11),
TO_SIGNED(373,11),
TO_SIGNED(331,11),
TO_SIGNED(288,11),
TO_SIGNED(244,11),
TO_SIGNED(200,11),
TO_SIGNED(154,11),
TO_SIGNED(108,11),
TO_SIGNED(61,11),
TO_SIGNED(14,11),
TO_SIGNED(-33,11),
TO_SIGNED(-80,11),
TO_SIGNED(-127,11),
TO_SIGNED(-173,11),
TO_SIGNED(-218,11),
TO_SIGNED(-263,11),
TO_SIGNED(-306,11),
TO_SIGNED(-348,11),
TO_SIGNED(-389,11),
TO_SIGNED(-429,11),
TO_SIGNED(-466,11),
TO_SIGNED(-502,11),
TO_SIGNED(-536,11),
TO_SIGNED(-568,11),
TO_SIGNED(-598,11),
TO_SIGNED(-625,11),
TO_SIGNED(-650,11),
TO_SIGNED(-672,11),
TO_SIGNED(-691,11),
TO_SIGNED(-708,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-686,11),
TO_SIGNED(-665,11),
TO_SIGNED(-642,11),
TO_SIGNED(-617,11),
TO_SIGNED(-589,11),
TO_SIGNED(-559,11),
TO_SIGNED(-526,11),
TO_SIGNED(-492,11),
TO_SIGNED(-455,11),
TO_SIGNED(-417,11),
TO_SIGNED(-377,11),
TO_SIGNED(-336,11),
TO_SIGNED(-293,11),
TO_SIGNED(-249,11),
TO_SIGNED(-205,11),
TO_SIGNED(-159,11),
TO_SIGNED(-113,11),
TO_SIGNED(-66,11),
TO_SIGNED(-19,11),
TO_SIGNED(28,11),
TO_SIGNED(75,11),
TO_SIGNED(121,11),
TO_SIGNED(167,11),
TO_SIGNED(213,11),
TO_SIGNED(258,11),
TO_SIGNED(301,11),
TO_SIGNED(344,11),
TO_SIGNED(385,11),
TO_SIGNED(424,11),
TO_SIGNED(462,11),
TO_SIGNED(498,11),
TO_SIGNED(532,11),
TO_SIGNED(564,11),
TO_SIGNED(594,11),
TO_SIGNED(622,11),
TO_SIGNED(647,11),
TO_SIGNED(669,11),
TO_SIGNED(689,11),
TO_SIGNED(706,11),
TO_SIGNED(721,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(720,11),
TO_SIGNED(705,11),
TO_SIGNED(688,11),
TO_SIGNED(668,11),
TO_SIGNED(645,11),
TO_SIGNED(620,11),
TO_SIGNED(592,11),
TO_SIGNED(562,11),
TO_SIGNED(530,11),
TO_SIGNED(496,11),
TO_SIGNED(460,11),
TO_SIGNED(422,11),
TO_SIGNED(382,11),
TO_SIGNED(341,11),
TO_SIGNED(298,11),
TO_SIGNED(255,11),
TO_SIGNED(210,11),
TO_SIGNED(164,11),
TO_SIGNED(118,11),
TO_SIGNED(71,11),
TO_SIGNED(25,11),
TO_SIGNED(-22,11),
TO_SIGNED(-69,11),
TO_SIGNED(-116,11),
TO_SIGNED(-162,11),
TO_SIGNED(-208,11),
TO_SIGNED(-252,11),
TO_SIGNED(-296,11),
TO_SIGNED(-339,11),
TO_SIGNED(-380,11),
TO_SIGNED(-420,11),
TO_SIGNED(-458,11),
TO_SIGNED(-494,11),
TO_SIGNED(-529,11),
TO_SIGNED(-561,11),
TO_SIGNED(-591,11),
TO_SIGNED(-619,11),
TO_SIGNED(-644,11),
TO_SIGNED(-667,11),
TO_SIGNED(-687,11),
TO_SIGNED(-705,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-733,11),
TO_SIGNED(-721,11),
TO_SIGNED(-707,11),
TO_SIGNED(-690,11),
TO_SIGNED(-670,11),
TO_SIGNED(-648,11),
TO_SIGNED(-623,11),
TO_SIGNED(-596,11),
TO_SIGNED(-566,11),
TO_SIGNED(-534,11),
TO_SIGNED(-500,11),
TO_SIGNED(-464,11),
TO_SIGNED(-426,11),
TO_SIGNED(-387,11),
TO_SIGNED(-345,11),
TO_SIGNED(-303,11),
TO_SIGNED(-260,11),
TO_SIGNED(-215,11),
TO_SIGNED(-169,11),
TO_SIGNED(-123,11),
TO_SIGNED(-77,11),
TO_SIGNED(-30,11),
TO_SIGNED(17,11),
TO_SIGNED(64,11),
TO_SIGNED(111,11),
TO_SIGNED(157,11),
TO_SIGNED(203,11),
TO_SIGNED(247,11),
TO_SIGNED(291,11),
TO_SIGNED(334,11),
TO_SIGNED(375,11),
TO_SIGNED(415,11),
TO_SIGNED(454,11),
TO_SIGNED(490,11),
TO_SIGNED(525,11),
TO_SIGNED(557,11),
TO_SIGNED(588,11),
TO_SIGNED(616,11),
TO_SIGNED(641,11),
TO_SIGNED(664,11),
TO_SIGNED(685,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(709,11),
TO_SIGNED(692,11),
TO_SIGNED(673,11),
TO_SIGNED(651,11),
TO_SIGNED(626,11),
TO_SIGNED(599,11),
TO_SIGNED(569,11),
TO_SIGNED(538,11),
TO_SIGNED(504,11),
TO_SIGNED(468,11),
TO_SIGNED(430,11),
TO_SIGNED(391,11),
TO_SIGNED(350,11),
TO_SIGNED(308,11),
TO_SIGNED(265,11),
TO_SIGNED(220,11),
TO_SIGNED(175,11),
TO_SIGNED(129,11),
TO_SIGNED(82,11),
TO_SIGNED(35,11),
TO_SIGNED(-12,11),
TO_SIGNED(-59,11),
TO_SIGNED(-105,11),
TO_SIGNED(-152,11),
TO_SIGNED(-197,11),
TO_SIGNED(-242,11),
TO_SIGNED(-286,11),
TO_SIGNED(-329,11),
TO_SIGNED(-371,11),
TO_SIGNED(-411,11),
TO_SIGNED(-449,11),
TO_SIGNED(-486,11),
TO_SIGNED(-521,11),
TO_SIGNED(-554,11),
TO_SIGNED(-584,11),
TO_SIGNED(-613,11),
TO_SIGNED(-639,11),
TO_SIGNED(-662,11),
TO_SIGNED(-683,11),
TO_SIGNED(-701,11),
TO_SIGNED(-716,11),
TO_SIGNED(-729,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-711,11),
TO_SIGNED(-694,11),
TO_SIGNED(-675,11),
TO_SIGNED(-653,11),
TO_SIGNED(-629,11),
TO_SIGNED(-602,11),
TO_SIGNED(-573,11),
TO_SIGNED(-541,11),
TO_SIGNED(-508,11),
TO_SIGNED(-472,11),
TO_SIGNED(-435,11),
TO_SIGNED(-396,11),
TO_SIGNED(-355,11),
TO_SIGNED(-313,11),
TO_SIGNED(-270,11),
TO_SIGNED(-225,11),
TO_SIGNED(-180,11),
TO_SIGNED(-134,11),
TO_SIGNED(-87,11),
TO_SIGNED(-41,11),
TO_SIGNED(6,11),
TO_SIGNED(53,11),
TO_SIGNED(100,11),
TO_SIGNED(147,11),
TO_SIGNED(192,11),
TO_SIGNED(237,11),
TO_SIGNED(281,11),
TO_SIGNED(324,11),
TO_SIGNED(366,11),
TO_SIGNED(406,11),
TO_SIGNED(445,11),
TO_SIGNED(482,11),
TO_SIGNED(517,11),
TO_SIGNED(550,11),
TO_SIGNED(581,11),
TO_SIGNED(610,11),
TO_SIGNED(636,11),
TO_SIGNED(659,11),
TO_SIGNED(681,11),
TO_SIGNED(699,11),
TO_SIGNED(715,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(712,11),
TO_SIGNED(696,11),
TO_SIGNED(677,11),
TO_SIGNED(656,11),
TO_SIGNED(632,11),
TO_SIGNED(605,11),
TO_SIGNED(576,11),
TO_SIGNED(545,11),
TO_SIGNED(512,11),
TO_SIGNED(476,11),
TO_SIGNED(439,11),
TO_SIGNED(400,11),
TO_SIGNED(360,11),
TO_SIGNED(318,11),
TO_SIGNED(275,11),
TO_SIGNED(230,11),
TO_SIGNED(185,11),
TO_SIGNED(139,11),
TO_SIGNED(93,11),
TO_SIGNED(46,11),
TO_SIGNED(-1,11),
TO_SIGNED(-48,11),
TO_SIGNED(-95,11),
TO_SIGNED(-141,11),
TO_SIGNED(-187,11),
TO_SIGNED(-232,11),
TO_SIGNED(-276,11),
TO_SIGNED(-320,11),
TO_SIGNED(-362,11),
TO_SIGNED(-402,11),
TO_SIGNED(-441,11),
TO_SIGNED(-478,11),
TO_SIGNED(-513,11),
TO_SIGNED(-547,11),
TO_SIGNED(-578,11),
TO_SIGNED(-606,11),
TO_SIGNED(-633,11),
TO_SIGNED(-657,11),
TO_SIGNED(-678,11),
TO_SIGNED(-697,11),
TO_SIGNED(-713,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-714,11),
TO_SIGNED(-698,11),
TO_SIGNED(-680,11),
TO_SIGNED(-658,11),
TO_SIGNED(-635,11),
TO_SIGNED(-608,11),
TO_SIGNED(-580,11),
TO_SIGNED(-549,11),
TO_SIGNED(-516,11),
TO_SIGNED(-480,11),
TO_SIGNED(-443,11),
TO_SIGNED(-405,11),
TO_SIGNED(-364,11),
TO_SIGNED(-323,11),
TO_SIGNED(-279,11),
TO_SIGNED(-235,11),
TO_SIGNED(-190,11),
TO_SIGNED(-144,11),
TO_SIGNED(-98,11),
TO_SIGNED(-51,11),
TO_SIGNED(-4,11),
TO_SIGNED(43,11),
TO_SIGNED(90,11),
TO_SIGNED(136,11),
TO_SIGNED(182,11),
TO_SIGNED(227,11),
TO_SIGNED(272,11),
TO_SIGNED(315,11),
TO_SIGNED(357,11),
TO_SIGNED(397,11),
TO_SIGNED(437,11),
TO_SIGNED(474,11),
TO_SIGNED(509,11),
TO_SIGNED(543,11),
TO_SIGNED(574,11),
TO_SIGNED(603,11),
TO_SIGNED(630,11),
TO_SIGNED(654,11),
TO_SIGNED(676,11),
TO_SIGNED(695,11),
TO_SIGNED(711,11),
TO_SIGNED(725,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(716,11),
TO_SIGNED(700,11),
TO_SIGNED(682,11),
TO_SIGNED(661,11),
TO_SIGNED(637,11),
TO_SIGNED(611,11),
TO_SIGNED(583,11),
TO_SIGNED(552,11),
TO_SIGNED(519,11),
TO_SIGNED(485,11),
TO_SIGNED(448,11),
TO_SIGNED(409,11),
TO_SIGNED(369,11),
TO_SIGNED(327,11),
TO_SIGNED(284,11),
TO_SIGNED(240,11),
TO_SIGNED(195,11),
TO_SIGNED(150,11),
TO_SIGNED(103,11),
TO_SIGNED(57,11),
TO_SIGNED(10,11),
TO_SIGNED(-37,11),
TO_SIGNED(-84,11),
TO_SIGNED(-131,11),
TO_SIGNED(-177,11),
TO_SIGNED(-222,11),
TO_SIGNED(-267,11),
TO_SIGNED(-310,11),
TO_SIGNED(-352,11),
TO_SIGNED(-393,11),
TO_SIGNED(-432,11),
TO_SIGNED(-470,11),
TO_SIGNED(-505,11),
TO_SIGNED(-539,11),
TO_SIGNED(-571,11),
TO_SIGNED(-600,11),
TO_SIGNED(-627,11),
TO_SIGNED(-652,11),
TO_SIGNED(-674,11),
TO_SIGNED(-693,11),
TO_SIGNED(-710,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-702,11),
TO_SIGNED(-684,11),
TO_SIGNED(-663,11),
TO_SIGNED(-640,11),
TO_SIGNED(-615,11),
TO_SIGNED(-586,11),
TO_SIGNED(-556,11),
TO_SIGNED(-523,11),
TO_SIGNED(-489,11),
TO_SIGNED(-452,11),
TO_SIGNED(-414,11),
TO_SIGNED(-374,11),
TO_SIGNED(-332,11),
TO_SIGNED(-289,11),
TO_SIGNED(-245,11),
TO_SIGNED(-201,11),
TO_SIGNED(-155,11),
TO_SIGNED(-109,11),
TO_SIGNED(-62,11),
TO_SIGNED(-15,11),
TO_SIGNED(32,11),
TO_SIGNED(79,11),
TO_SIGNED(125,11),
TO_SIGNED(172,11),
TO_SIGNED(217,11),
TO_SIGNED(262,11),
TO_SIGNED(305,11),
TO_SIGNED(347,11),
TO_SIGNED(388,11),
TO_SIGNED(428,11),
TO_SIGNED(466,11),
TO_SIGNED(501,11),
TO_SIGNED(535,11),
TO_SIGNED(567,11),
TO_SIGNED(597,11),
TO_SIGNED(624,11),
TO_SIGNED(649,11),
TO_SIGNED(671,11),
TO_SIGNED(691,11),
TO_SIGNED(708,11),
TO_SIGNED(722,11),
TO_SIGNED(733,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(704,11),
TO_SIGNED(686,11),
TO_SIGNED(666,11),
TO_SIGNED(643,11),
TO_SIGNED(618,11),
TO_SIGNED(590,11),
TO_SIGNED(559,11),
TO_SIGNED(527,11),
TO_SIGNED(493,11),
TO_SIGNED(456,11),
TO_SIGNED(418,11),
TO_SIGNED(378,11),
TO_SIGNED(337,11),
TO_SIGNED(294,11),
TO_SIGNED(250,11),
TO_SIGNED(206,11),
TO_SIGNED(160,11),
TO_SIGNED(114,11),
TO_SIGNED(67,11),
TO_SIGNED(20,11),
TO_SIGNED(-27,11),
TO_SIGNED(-74,11),
TO_SIGNED(-120,11),
TO_SIGNED(-166,11),
TO_SIGNED(-212,11),
TO_SIGNED(-257,11),
TO_SIGNED(-300,11),
TO_SIGNED(-343,11),
TO_SIGNED(-384,11),
TO_SIGNED(-423,11),
TO_SIGNED(-461,11),
TO_SIGNED(-497,11),
TO_SIGNED(-532,11),
TO_SIGNED(-564,11),
TO_SIGNED(-594,11),
TO_SIGNED(-621,11),
TO_SIGNED(-646,11),
TO_SIGNED(-669,11),
TO_SIGNED(-689,11),
TO_SIGNED(-706,11),
TO_SIGNED(-721,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-720,11),
TO_SIGNED(-706,11),
TO_SIGNED(-688,11),
TO_SIGNED(-668,11),
TO_SIGNED(-646,11),
TO_SIGNED(-621,11),
TO_SIGNED(-593,11),
TO_SIGNED(-563,11),
TO_SIGNED(-531,11),
TO_SIGNED(-497,11),
TO_SIGNED(-460,11),
TO_SIGNED(-422,11),
TO_SIGNED(-383,11),
TO_SIGNED(-342,11),
TO_SIGNED(-299,11),
TO_SIGNED(-256,11),
TO_SIGNED(-211,11),
TO_SIGNED(-165,11),
TO_SIGNED(-119,11),
TO_SIGNED(-73,11),
TO_SIGNED(-26,11),
TO_SIGNED(21,11),
TO_SIGNED(68,11),
TO_SIGNED(115,11),
TO_SIGNED(161,11),
TO_SIGNED(207,11),
TO_SIGNED(251,11),
TO_SIGNED(295,11),
TO_SIGNED(338,11),
TO_SIGNED(379,11),
TO_SIGNED(419,11),
TO_SIGNED(457,11),
TO_SIGNED(493,11),
TO_SIGNED(528,11),
TO_SIGNED(560,11),
TO_SIGNED(590,11),
TO_SIGNED(618,11),
TO_SIGNED(644,11),
TO_SIGNED(666,11),
TO_SIGNED(687,11),
TO_SIGNED(704,11),
TO_SIGNED(719,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(671,11),
TO_SIGNED(648,11),
TO_SIGNED(624,11),
TO_SIGNED(596,11),
TO_SIGNED(567,11),
TO_SIGNED(535,11),
TO_SIGNED(501,11),
TO_SIGNED(465,11),
TO_SIGNED(427,11),
TO_SIGNED(387,11),
TO_SIGNED(346,11),
TO_SIGNED(304,11),
TO_SIGNED(261,11),
TO_SIGNED(216,11),
TO_SIGNED(171,11),
TO_SIGNED(124,11),
TO_SIGNED(78,11),
TO_SIGNED(31,11),
TO_SIGNED(-16,11),
TO_SIGNED(-63,11),
TO_SIGNED(-110,11),
TO_SIGNED(-156,11),
TO_SIGNED(-202,11),
TO_SIGNED(-246,11),
TO_SIGNED(-290,11),
TO_SIGNED(-333,11),
TO_SIGNED(-375,11),
TO_SIGNED(-415,11),
TO_SIGNED(-453,11),
TO_SIGNED(-489,11),
TO_SIGNED(-524,11),
TO_SIGNED(-557,11),
TO_SIGNED(-587,11),
TO_SIGNED(-615,11),
TO_SIGNED(-641,11),
TO_SIGNED(-664,11),
TO_SIGNED(-685,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-730,11),
TO_SIGNED(-739,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-693,11),
TO_SIGNED(-673,11),
TO_SIGNED(-651,11),
TO_SIGNED(-627,11),
TO_SIGNED(-599,11),
TO_SIGNED(-570,11),
TO_SIGNED(-538,11),
TO_SIGNED(-505,11),
TO_SIGNED(-469,11),
TO_SIGNED(-431,11),
TO_SIGNED(-392,11),
TO_SIGNED(-351,11),
TO_SIGNED(-309,11),
TO_SIGNED(-266,11),
TO_SIGNED(-221,11),
TO_SIGNED(-176,11),
TO_SIGNED(-130,11),
TO_SIGNED(-83,11),
TO_SIGNED(-36,11),
TO_SIGNED(11,11),
TO_SIGNED(58,11),
TO_SIGNED(104,11),
TO_SIGNED(151,11),
TO_SIGNED(196,11),
TO_SIGNED(241,11),
TO_SIGNED(285,11),
TO_SIGNED(328,11),
TO_SIGNED(370,11),
TO_SIGNED(410,11),
TO_SIGNED(449,11),
TO_SIGNED(485,11),
TO_SIGNED(520,11),
TO_SIGNED(553,11),
TO_SIGNED(584,11),
TO_SIGNED(612,11),
TO_SIGNED(638,11),
TO_SIGNED(661,11),
TO_SIGNED(682,11),
TO_SIGNED(700,11),
TO_SIGNED(716,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(725,11),
TO_SIGNED(711,11),
TO_SIGNED(695,11),
TO_SIGNED(675,11),
TO_SIGNED(654,11),
TO_SIGNED(629,11),
TO_SIGNED(603,11),
TO_SIGNED(574,11),
TO_SIGNED(542,11),
TO_SIGNED(509,11),
TO_SIGNED(473,11),
TO_SIGNED(436,11),
TO_SIGNED(397,11),
TO_SIGNED(356,11),
TO_SIGNED(314,11),
TO_SIGNED(271,11),
TO_SIGNED(226,11),
TO_SIGNED(181,11),
TO_SIGNED(135,11),
TO_SIGNED(88,11),
TO_SIGNED(42,11),
TO_SIGNED(-5,11),
TO_SIGNED(-52,11),
TO_SIGNED(-99,11),
TO_SIGNED(-145,11),
TO_SIGNED(-191,11),
TO_SIGNED(-236,11),
TO_SIGNED(-280,11),
TO_SIGNED(-323,11),
TO_SIGNED(-365,11),
TO_SIGNED(-406,11),
TO_SIGNED(-444,11),
TO_SIGNED(-481,11),
TO_SIGNED(-516,11),
TO_SIGNED(-549,11),
TO_SIGNED(-580,11),
TO_SIGNED(-609,11),
TO_SIGNED(-635,11),
TO_SIGNED(-659,11),
TO_SIGNED(-680,11),
TO_SIGNED(-699,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-736,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-678,11),
TO_SIGNED(-656,11),
TO_SIGNED(-632,11),
TO_SIGNED(-606,11),
TO_SIGNED(-577,11),
TO_SIGNED(-546,11),
TO_SIGNED(-512,11),
TO_SIGNED(-477,11),
TO_SIGNED(-440,11),
TO_SIGNED(-401,11),
TO_SIGNED(-361,11),
TO_SIGNED(-319,11),
TO_SIGNED(-275,11),
TO_SIGNED(-231,11),
TO_SIGNED(-186,11),
TO_SIGNED(-140,11),
TO_SIGNED(-94,11),
TO_SIGNED(-47,11),
TO_SIGNED(0,11),
TO_SIGNED(47,11),
TO_SIGNED(94,11),
TO_SIGNED(140,11),
TO_SIGNED(186,11),
TO_SIGNED(231,11),
TO_SIGNED(275,11),
TO_SIGNED(319,11),
TO_SIGNED(361,11),
TO_SIGNED(401,11),
TO_SIGNED(440,11),
TO_SIGNED(477,11),
TO_SIGNED(512,11),
TO_SIGNED(546,11),
TO_SIGNED(577,11),
TO_SIGNED(606,11),
TO_SIGNED(632,11),
TO_SIGNED(656,11),
TO_SIGNED(678,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(736,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(699,11),
TO_SIGNED(680,11),
TO_SIGNED(659,11),
TO_SIGNED(635,11),
TO_SIGNED(609,11),
TO_SIGNED(580,11),
TO_SIGNED(549,11),
TO_SIGNED(516,11),
TO_SIGNED(481,11),
TO_SIGNED(444,11),
TO_SIGNED(406,11),
TO_SIGNED(365,11),
TO_SIGNED(323,11),
TO_SIGNED(280,11),
TO_SIGNED(236,11),
TO_SIGNED(191,11),
TO_SIGNED(145,11),
TO_SIGNED(99,11),
TO_SIGNED(52,11),
TO_SIGNED(5,11),
TO_SIGNED(-42,11),
TO_SIGNED(-88,11),
TO_SIGNED(-135,11),
TO_SIGNED(-181,11),
TO_SIGNED(-226,11),
TO_SIGNED(-271,11),
TO_SIGNED(-314,11),
TO_SIGNED(-356,11),
TO_SIGNED(-397,11),
TO_SIGNED(-436,11),
TO_SIGNED(-473,11),
TO_SIGNED(-509,11),
TO_SIGNED(-542,11),
TO_SIGNED(-574,11),
TO_SIGNED(-603,11),
TO_SIGNED(-629,11),
TO_SIGNED(-654,11),
TO_SIGNED(-675,11),
TO_SIGNED(-695,11),
TO_SIGNED(-711,11),
TO_SIGNED(-725,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-716,11),
TO_SIGNED(-700,11),
TO_SIGNED(-682,11),
TO_SIGNED(-661,11),
TO_SIGNED(-638,11),
TO_SIGNED(-612,11),
TO_SIGNED(-584,11),
TO_SIGNED(-553,11),
TO_SIGNED(-520,11),
TO_SIGNED(-485,11),
TO_SIGNED(-449,11),
TO_SIGNED(-410,11),
TO_SIGNED(-370,11),
TO_SIGNED(-328,11),
TO_SIGNED(-285,11),
TO_SIGNED(-241,11),
TO_SIGNED(-196,11),
TO_SIGNED(-151,11),
TO_SIGNED(-104,11),
TO_SIGNED(-58,11),
TO_SIGNED(-11,11),
TO_SIGNED(36,11),
TO_SIGNED(83,11),
TO_SIGNED(130,11),
TO_SIGNED(176,11),
TO_SIGNED(221,11),
TO_SIGNED(266,11),
TO_SIGNED(309,11),
TO_SIGNED(351,11),
TO_SIGNED(392,11),
TO_SIGNED(431,11),
TO_SIGNED(469,11),
TO_SIGNED(505,11),
TO_SIGNED(538,11),
TO_SIGNED(570,11),
TO_SIGNED(599,11),
TO_SIGNED(627,11),
TO_SIGNED(651,11),
TO_SIGNED(673,11),
TO_SIGNED(693,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(739,11),
TO_SIGNED(730,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(685,11),
TO_SIGNED(664,11),
TO_SIGNED(641,11),
TO_SIGNED(615,11),
TO_SIGNED(587,11),
TO_SIGNED(557,11),
TO_SIGNED(524,11),
TO_SIGNED(489,11),
TO_SIGNED(453,11),
TO_SIGNED(415,11),
TO_SIGNED(375,11),
TO_SIGNED(333,11),
TO_SIGNED(290,11),
TO_SIGNED(246,11),
TO_SIGNED(202,11),
TO_SIGNED(156,11),
TO_SIGNED(110,11),
TO_SIGNED(63,11),
TO_SIGNED(16,11),
TO_SIGNED(-31,11),
TO_SIGNED(-78,11),
TO_SIGNED(-124,11),
TO_SIGNED(-171,11),
TO_SIGNED(-216,11),
TO_SIGNED(-261,11),
TO_SIGNED(-304,11),
TO_SIGNED(-346,11),
TO_SIGNED(-387,11),
TO_SIGNED(-427,11),
TO_SIGNED(-465,11),
TO_SIGNED(-501,11),
TO_SIGNED(-535,11),
TO_SIGNED(-567,11),
TO_SIGNED(-596,11),
TO_SIGNED(-624,11),
TO_SIGNED(-648,11),
TO_SIGNED(-671,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-719,11),
TO_SIGNED(-704,11),
TO_SIGNED(-687,11),
TO_SIGNED(-666,11),
TO_SIGNED(-644,11),
TO_SIGNED(-618,11),
TO_SIGNED(-590,11),
TO_SIGNED(-560,11),
TO_SIGNED(-528,11),
TO_SIGNED(-493,11),
TO_SIGNED(-457,11),
TO_SIGNED(-419,11),
TO_SIGNED(-379,11),
TO_SIGNED(-338,11),
TO_SIGNED(-295,11),
TO_SIGNED(-251,11),
TO_SIGNED(-207,11),
TO_SIGNED(-161,11),
TO_SIGNED(-115,11),
TO_SIGNED(-68,11),
TO_SIGNED(-21,11),
TO_SIGNED(26,11),
TO_SIGNED(73,11),
TO_SIGNED(119,11),
TO_SIGNED(165,11),
TO_SIGNED(211,11),
TO_SIGNED(256,11),
TO_SIGNED(299,11),
TO_SIGNED(342,11),
TO_SIGNED(383,11),
TO_SIGNED(422,11),
TO_SIGNED(460,11),
TO_SIGNED(497,11),
TO_SIGNED(531,11),
TO_SIGNED(563,11),
TO_SIGNED(593,11),
TO_SIGNED(621,11),
TO_SIGNED(646,11),
TO_SIGNED(668,11),
TO_SIGNED(688,11),
TO_SIGNED(706,11),
TO_SIGNED(720,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(721,11),
TO_SIGNED(706,11),
TO_SIGNED(689,11),
TO_SIGNED(669,11),
TO_SIGNED(646,11),
TO_SIGNED(621,11),
TO_SIGNED(594,11),
TO_SIGNED(564,11),
TO_SIGNED(532,11),
TO_SIGNED(497,11),
TO_SIGNED(461,11),
TO_SIGNED(423,11),
TO_SIGNED(384,11),
TO_SIGNED(343,11),
TO_SIGNED(300,11),
TO_SIGNED(257,11),
TO_SIGNED(212,11),
TO_SIGNED(166,11),
TO_SIGNED(120,11),
TO_SIGNED(74,11),
TO_SIGNED(27,11),
TO_SIGNED(-20,11),
TO_SIGNED(-67,11),
TO_SIGNED(-114,11),
TO_SIGNED(-160,11),
TO_SIGNED(-206,11),
TO_SIGNED(-250,11),
TO_SIGNED(-294,11),
TO_SIGNED(-337,11),
TO_SIGNED(-378,11),
TO_SIGNED(-418,11),
TO_SIGNED(-456,11),
TO_SIGNED(-493,11),
TO_SIGNED(-527,11),
TO_SIGNED(-559,11),
TO_SIGNED(-590,11),
TO_SIGNED(-618,11),
TO_SIGNED(-643,11),
TO_SIGNED(-666,11),
TO_SIGNED(-686,11),
TO_SIGNED(-704,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-733,11),
TO_SIGNED(-722,11),
TO_SIGNED(-708,11),
TO_SIGNED(-691,11),
TO_SIGNED(-671,11),
TO_SIGNED(-649,11),
TO_SIGNED(-624,11),
TO_SIGNED(-597,11),
TO_SIGNED(-567,11),
TO_SIGNED(-535,11),
TO_SIGNED(-501,11),
TO_SIGNED(-466,11),
TO_SIGNED(-428,11),
TO_SIGNED(-388,11),
TO_SIGNED(-347,11),
TO_SIGNED(-305,11),
TO_SIGNED(-262,11),
TO_SIGNED(-217,11),
TO_SIGNED(-172,11),
TO_SIGNED(-125,11),
TO_SIGNED(-79,11),
TO_SIGNED(-32,11),
TO_SIGNED(15,11),
TO_SIGNED(62,11),
TO_SIGNED(109,11),
TO_SIGNED(155,11),
TO_SIGNED(201,11),
TO_SIGNED(245,11),
TO_SIGNED(289,11),
TO_SIGNED(332,11),
TO_SIGNED(374,11),
TO_SIGNED(414,11),
TO_SIGNED(452,11),
TO_SIGNED(489,11),
TO_SIGNED(523,11),
TO_SIGNED(556,11),
TO_SIGNED(586,11),
TO_SIGNED(615,11),
TO_SIGNED(640,11),
TO_SIGNED(663,11),
TO_SIGNED(684,11),
TO_SIGNED(702,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(710,11),
TO_SIGNED(693,11),
TO_SIGNED(674,11),
TO_SIGNED(652,11),
TO_SIGNED(627,11),
TO_SIGNED(600,11),
TO_SIGNED(571,11),
TO_SIGNED(539,11),
TO_SIGNED(505,11),
TO_SIGNED(470,11),
TO_SIGNED(432,11),
TO_SIGNED(393,11),
TO_SIGNED(352,11),
TO_SIGNED(310,11),
TO_SIGNED(267,11),
TO_SIGNED(222,11),
TO_SIGNED(177,11),
TO_SIGNED(131,11),
TO_SIGNED(84,11),
TO_SIGNED(37,11),
TO_SIGNED(-10,11),
TO_SIGNED(-57,11),
TO_SIGNED(-103,11),
TO_SIGNED(-150,11),
TO_SIGNED(-195,11),
TO_SIGNED(-240,11),
TO_SIGNED(-284,11),
TO_SIGNED(-327,11),
TO_SIGNED(-369,11),
TO_SIGNED(-409,11),
TO_SIGNED(-448,11),
TO_SIGNED(-485,11),
TO_SIGNED(-519,11),
TO_SIGNED(-552,11),
TO_SIGNED(-583,11),
TO_SIGNED(-611,11),
TO_SIGNED(-637,11),
TO_SIGNED(-661,11),
TO_SIGNED(-682,11),
TO_SIGNED(-700,11),
TO_SIGNED(-716,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-725,11),
TO_SIGNED(-711,11),
TO_SIGNED(-695,11),
TO_SIGNED(-676,11),
TO_SIGNED(-654,11),
TO_SIGNED(-630,11),
TO_SIGNED(-603,11),
TO_SIGNED(-574,11),
TO_SIGNED(-543,11),
TO_SIGNED(-509,11),
TO_SIGNED(-474,11),
TO_SIGNED(-437,11),
TO_SIGNED(-397,11),
TO_SIGNED(-357,11),
TO_SIGNED(-315,11),
TO_SIGNED(-272,11),
TO_SIGNED(-227,11),
TO_SIGNED(-182,11),
TO_SIGNED(-136,11),
TO_SIGNED(-90,11),
TO_SIGNED(-43,11),
TO_SIGNED(4,11),
TO_SIGNED(51,11),
TO_SIGNED(98,11),
TO_SIGNED(144,11),
TO_SIGNED(190,11),
TO_SIGNED(235,11),
TO_SIGNED(279,11),
TO_SIGNED(323,11),
TO_SIGNED(364,11),
TO_SIGNED(405,11),
TO_SIGNED(443,11),
TO_SIGNED(480,11),
TO_SIGNED(516,11),
TO_SIGNED(549,11),
TO_SIGNED(580,11),
TO_SIGNED(608,11),
TO_SIGNED(635,11),
TO_SIGNED(658,11),
TO_SIGNED(680,11),
TO_SIGNED(698,11),
TO_SIGNED(714,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(713,11),
TO_SIGNED(697,11),
TO_SIGNED(678,11),
TO_SIGNED(657,11),
TO_SIGNED(633,11),
TO_SIGNED(606,11),
TO_SIGNED(578,11),
TO_SIGNED(547,11),
TO_SIGNED(513,11),
TO_SIGNED(478,11),
TO_SIGNED(441,11),
TO_SIGNED(402,11),
TO_SIGNED(362,11),
TO_SIGNED(320,11),
TO_SIGNED(276,11),
TO_SIGNED(232,11),
TO_SIGNED(187,11),
TO_SIGNED(141,11),
TO_SIGNED(95,11),
TO_SIGNED(48,11),
TO_SIGNED(1,11),
TO_SIGNED(-46,11),
TO_SIGNED(-93,11),
TO_SIGNED(-139,11),
TO_SIGNED(-185,11),
TO_SIGNED(-230,11),
TO_SIGNED(-275,11),
TO_SIGNED(-318,11),
TO_SIGNED(-360,11),
TO_SIGNED(-400,11),
TO_SIGNED(-439,11),
TO_SIGNED(-476,11),
TO_SIGNED(-512,11),
TO_SIGNED(-545,11),
TO_SIGNED(-576,11),
TO_SIGNED(-605,11),
TO_SIGNED(-632,11),
TO_SIGNED(-656,11),
TO_SIGNED(-677,11),
TO_SIGNED(-696,11),
TO_SIGNED(-712,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-715,11),
TO_SIGNED(-699,11),
TO_SIGNED(-681,11),
TO_SIGNED(-659,11),
TO_SIGNED(-636,11),
TO_SIGNED(-610,11),
TO_SIGNED(-581,11),
TO_SIGNED(-550,11),
TO_SIGNED(-517,11),
TO_SIGNED(-482,11),
TO_SIGNED(-445,11),
TO_SIGNED(-406,11),
TO_SIGNED(-366,11),
TO_SIGNED(-324,11),
TO_SIGNED(-281,11),
TO_SIGNED(-237,11),
TO_SIGNED(-192,11),
TO_SIGNED(-147,11),
TO_SIGNED(-100,11),
TO_SIGNED(-53,11),
TO_SIGNED(-6,11),
TO_SIGNED(41,11),
TO_SIGNED(87,11),
TO_SIGNED(134,11),
TO_SIGNED(180,11),
TO_SIGNED(225,11),
TO_SIGNED(270,11),
TO_SIGNED(313,11),
TO_SIGNED(355,11),
TO_SIGNED(396,11),
TO_SIGNED(435,11),
TO_SIGNED(472,11),
TO_SIGNED(508,11),
TO_SIGNED(541,11),
TO_SIGNED(573,11),
TO_SIGNED(602,11),
TO_SIGNED(629,11),
TO_SIGNED(653,11),
TO_SIGNED(675,11),
TO_SIGNED(694,11),
TO_SIGNED(711,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(729,11),
TO_SIGNED(716,11),
TO_SIGNED(701,11),
TO_SIGNED(683,11),
TO_SIGNED(662,11),
TO_SIGNED(639,11),
TO_SIGNED(613,11),
TO_SIGNED(584,11),
TO_SIGNED(554,11),
TO_SIGNED(521,11),
TO_SIGNED(486,11),
TO_SIGNED(449,11),
TO_SIGNED(411,11),
TO_SIGNED(371,11),
TO_SIGNED(329,11),
TO_SIGNED(286,11),
TO_SIGNED(242,11),
TO_SIGNED(197,11),
TO_SIGNED(152,11),
TO_SIGNED(105,11),
TO_SIGNED(59,11),
TO_SIGNED(12,11),
TO_SIGNED(-35,11),
TO_SIGNED(-82,11),
TO_SIGNED(-129,11),
TO_SIGNED(-175,11),
TO_SIGNED(-220,11),
TO_SIGNED(-265,11),
TO_SIGNED(-308,11),
TO_SIGNED(-350,11),
TO_SIGNED(-391,11),
TO_SIGNED(-430,11),
TO_SIGNED(-468,11),
TO_SIGNED(-504,11),
TO_SIGNED(-538,11),
TO_SIGNED(-569,11),
TO_SIGNED(-599,11),
TO_SIGNED(-626,11),
TO_SIGNED(-651,11),
TO_SIGNED(-673,11),
TO_SIGNED(-692,11),
TO_SIGNED(-709,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-685,11),
TO_SIGNED(-664,11),
TO_SIGNED(-641,11),
TO_SIGNED(-616,11),
TO_SIGNED(-588,11),
TO_SIGNED(-557,11),
TO_SIGNED(-525,11),
TO_SIGNED(-490,11),
TO_SIGNED(-454,11),
TO_SIGNED(-415,11),
TO_SIGNED(-375,11),
TO_SIGNED(-334,11),
TO_SIGNED(-291,11),
TO_SIGNED(-247,11),
TO_SIGNED(-203,11),
TO_SIGNED(-157,11),
TO_SIGNED(-111,11),
TO_SIGNED(-64,11),
TO_SIGNED(-17,11),
TO_SIGNED(30,11),
TO_SIGNED(77,11),
TO_SIGNED(123,11),
TO_SIGNED(169,11),
TO_SIGNED(215,11),
TO_SIGNED(260,11),
TO_SIGNED(303,11),
TO_SIGNED(345,11),
TO_SIGNED(387,11),
TO_SIGNED(426,11),
TO_SIGNED(464,11),
TO_SIGNED(500,11),
TO_SIGNED(534,11),
TO_SIGNED(566,11),
TO_SIGNED(596,11),
TO_SIGNED(623,11),
TO_SIGNED(648,11),
TO_SIGNED(670,11),
TO_SIGNED(690,11),
TO_SIGNED(707,11),
TO_SIGNED(721,11),
TO_SIGNED(733,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(705,11),
TO_SIGNED(687,11),
TO_SIGNED(667,11),
TO_SIGNED(644,11),
TO_SIGNED(619,11),
TO_SIGNED(591,11),
TO_SIGNED(561,11),
TO_SIGNED(529,11),
TO_SIGNED(494,11),
TO_SIGNED(458,11),
TO_SIGNED(420,11),
TO_SIGNED(380,11),
TO_SIGNED(339,11),
TO_SIGNED(296,11),
TO_SIGNED(252,11),
TO_SIGNED(208,11),
TO_SIGNED(162,11),
TO_SIGNED(116,11),
TO_SIGNED(69,11),
TO_SIGNED(22,11),
TO_SIGNED(-25,11),
TO_SIGNED(-71,11),
TO_SIGNED(-118,11),
TO_SIGNED(-164,11),
TO_SIGNED(-210,11),
TO_SIGNED(-255,11),
TO_SIGNED(-298,11),
TO_SIGNED(-341,11),
TO_SIGNED(-382,11),
TO_SIGNED(-422,11),
TO_SIGNED(-460,11),
TO_SIGNED(-496,11),
TO_SIGNED(-530,11),
TO_SIGNED(-562,11),
TO_SIGNED(-592,11),
TO_SIGNED(-620,11),
TO_SIGNED(-645,11),
TO_SIGNED(-668,11),
TO_SIGNED(-688,11),
TO_SIGNED(-705,11),
TO_SIGNED(-720,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-721,11),
TO_SIGNED(-706,11),
TO_SIGNED(-689,11),
TO_SIGNED(-669,11),
TO_SIGNED(-647,11),
TO_SIGNED(-622,11),
TO_SIGNED(-594,11),
TO_SIGNED(-564,11),
TO_SIGNED(-532,11),
TO_SIGNED(-498,11),
TO_SIGNED(-462,11),
TO_SIGNED(-424,11),
TO_SIGNED(-385,11),
TO_SIGNED(-344,11),
TO_SIGNED(-301,11),
TO_SIGNED(-258,11),
TO_SIGNED(-213,11),
TO_SIGNED(-167,11),
TO_SIGNED(-121,11),
TO_SIGNED(-75,11),
TO_SIGNED(-28,11),
TO_SIGNED(19,11),
TO_SIGNED(66,11),
TO_SIGNED(113,11),
TO_SIGNED(159,11),
TO_SIGNED(205,11),
TO_SIGNED(249,11),
TO_SIGNED(293,11),
TO_SIGNED(336,11),
TO_SIGNED(377,11),
TO_SIGNED(417,11),
TO_SIGNED(455,11),
TO_SIGNED(492,11),
TO_SIGNED(526,11),
TO_SIGNED(559,11),
TO_SIGNED(589,11),
TO_SIGNED(617,11),
TO_SIGNED(642,11),
TO_SIGNED(665,11),
TO_SIGNED(686,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(708,11),
TO_SIGNED(691,11),
TO_SIGNED(672,11),
TO_SIGNED(650,11),
TO_SIGNED(625,11),
TO_SIGNED(598,11),
TO_SIGNED(568,11),
TO_SIGNED(536,11),
TO_SIGNED(502,11),
TO_SIGNED(466,11),
TO_SIGNED(429,11),
TO_SIGNED(389,11),
TO_SIGNED(348,11),
TO_SIGNED(306,11),
TO_SIGNED(263,11),
TO_SIGNED(218,11),
TO_SIGNED(173,11),
TO_SIGNED(127,11),
TO_SIGNED(80,11),
TO_SIGNED(33,11),
TO_SIGNED(-14,11),
TO_SIGNED(-61,11),
TO_SIGNED(-108,11),
TO_SIGNED(-154,11),
TO_SIGNED(-200,11),
TO_SIGNED(-244,11),
TO_SIGNED(-288,11),
TO_SIGNED(-331,11),
TO_SIGNED(-373,11),
TO_SIGNED(-413,11),
TO_SIGNED(-451,11),
TO_SIGNED(-488,11),
TO_SIGNED(-523,11),
TO_SIGNED(-555,11),
TO_SIGNED(-586,11),
TO_SIGNED(-614,11),
TO_SIGNED(-640,11),
TO_SIGNED(-663,11),
TO_SIGNED(-684,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-729,11),
TO_SIGNED(-739,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-710,11),
TO_SIGNED(-693,11),
TO_SIGNED(-674,11),
TO_SIGNED(-652,11),
TO_SIGNED(-628,11),
TO_SIGNED(-601,11),
TO_SIGNED(-571,11),
TO_SIGNED(-540,11),
TO_SIGNED(-506,11),
TO_SIGNED(-471,11),
TO_SIGNED(-433,11),
TO_SIGNED(-394,11),
TO_SIGNED(-353,11),
TO_SIGNED(-311,11),
TO_SIGNED(-268,11),
TO_SIGNED(-223,11),
TO_SIGNED(-178,11),
TO_SIGNED(-132,11),
TO_SIGNED(-85,11),
TO_SIGNED(-38,11),
TO_SIGNED(9,11),
TO_SIGNED(56,11),
TO_SIGNED(102,11),
TO_SIGNED(149,11),
TO_SIGNED(194,11),
TO_SIGNED(239,11),
TO_SIGNED(283,11),
TO_SIGNED(326,11),
TO_SIGNED(368,11),
TO_SIGNED(408,11),
TO_SIGNED(447,11),
TO_SIGNED(484,11),
TO_SIGNED(519,11),
TO_SIGNED(552,11),
TO_SIGNED(582,11),
TO_SIGNED(611,11),
TO_SIGNED(637,11),
TO_SIGNED(660,11),
TO_SIGNED(681,11),
TO_SIGNED(700,11),
TO_SIGNED(715,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(736,11),
TO_SIGNED(725,11),
TO_SIGNED(712,11),
TO_SIGNED(695,11),
TO_SIGNED(676,11),
TO_SIGNED(655,11),
TO_SIGNED(631,11),
TO_SIGNED(604,11),
TO_SIGNED(575,11),
TO_SIGNED(544,11),
TO_SIGNED(510,11),
TO_SIGNED(475,11),
TO_SIGNED(437,11),
TO_SIGNED(398,11),
TO_SIGNED(358,11),
TO_SIGNED(316,11),
TO_SIGNED(273,11),
TO_SIGNED(228,11),
TO_SIGNED(183,11),
TO_SIGNED(137,11),
TO_SIGNED(91,11),
TO_SIGNED(44,11),
TO_SIGNED(-3,11),
TO_SIGNED(-50,11),
TO_SIGNED(-97,11),
TO_SIGNED(-143,11),
TO_SIGNED(-189,11),
TO_SIGNED(-234,11),
TO_SIGNED(-278,11),
TO_SIGNED(-322,11),
TO_SIGNED(-363,11),
TO_SIGNED(-404,11),
TO_SIGNED(-443,11),
TO_SIGNED(-480,11),
TO_SIGNED(-515,11),
TO_SIGNED(-548,11),
TO_SIGNED(-579,11),
TO_SIGNED(-608,11),
TO_SIGNED(-634,11),
TO_SIGNED(-658,11),
TO_SIGNED(-679,11),
TO_SIGNED(-698,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-679,11),
TO_SIGNED(-657,11),
TO_SIGNED(-633,11),
TO_SIGNED(-607,11),
TO_SIGNED(-578,11),
TO_SIGNED(-547,11),
TO_SIGNED(-514,11),
TO_SIGNED(-479,11),
TO_SIGNED(-442,11),
TO_SIGNED(-403,11),
TO_SIGNED(-362,11),
TO_SIGNED(-321,11),
TO_SIGNED(-277,11),
TO_SIGNED(-233,11),
TO_SIGNED(-188,11),
TO_SIGNED(-142,11),
TO_SIGNED(-96,11),
TO_SIGNED(-49,11),
TO_SIGNED(-2,11),
TO_SIGNED(45,11),
TO_SIGNED(92,11),
TO_SIGNED(138,11),
TO_SIGNED(184,11),
TO_SIGNED(229,11),
TO_SIGNED(274,11),
TO_SIGNED(317,11),
TO_SIGNED(359,11),
TO_SIGNED(399,11),
TO_SIGNED(438,11),
TO_SIGNED(476,11),
TO_SIGNED(511,11),
TO_SIGNED(544,11),
TO_SIGNED(576,11),
TO_SIGNED(605,11),
TO_SIGNED(631,11),
TO_SIGNED(655,11),
TO_SIGNED(677,11),
TO_SIGNED(696,11),
TO_SIGNED(712,11),
TO_SIGNED(725,11),
TO_SIGNED(736,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(715,11),
TO_SIGNED(699,11),
TO_SIGNED(681,11),
TO_SIGNED(660,11),
TO_SIGNED(636,11),
TO_SIGNED(610,11),
TO_SIGNED(582,11),
TO_SIGNED(551,11),
TO_SIGNED(518,11),
TO_SIGNED(483,11),
TO_SIGNED(446,11),
TO_SIGNED(407,11),
TO_SIGNED(367,11),
TO_SIGNED(325,11),
TO_SIGNED(282,11),
TO_SIGNED(238,11),
TO_SIGNED(193,11),
TO_SIGNED(148,11),
TO_SIGNED(101,11),
TO_SIGNED(54,11),
TO_SIGNED(7,11),
TO_SIGNED(-40,11),
TO_SIGNED(-86,11),
TO_SIGNED(-133,11),
TO_SIGNED(-179,11),
TO_SIGNED(-224,11),
TO_SIGNED(-269,11),
TO_SIGNED(-312,11),
TO_SIGNED(-354,11),
TO_SIGNED(-395,11),
TO_SIGNED(-434,11),
TO_SIGNED(-471,11),
TO_SIGNED(-507,11),
TO_SIGNED(-541,11),
TO_SIGNED(-572,11),
TO_SIGNED(-601,11),
TO_SIGNED(-628,11),
TO_SIGNED(-653,11),
TO_SIGNED(-675,11),
TO_SIGNED(-694,11),
TO_SIGNED(-710,11),
TO_SIGNED(-724,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-701,11),
TO_SIGNED(-683,11),
TO_SIGNED(-662,11),
TO_SIGNED(-639,11),
TO_SIGNED(-613,11),
TO_SIGNED(-585,11),
TO_SIGNED(-554,11),
TO_SIGNED(-522,11),
TO_SIGNED(-487,11),
TO_SIGNED(-450,11),
TO_SIGNED(-412,11),
TO_SIGNED(-372,11),
TO_SIGNED(-330,11),
TO_SIGNED(-287,11),
TO_SIGNED(-243,11),
TO_SIGNED(-198,11),
TO_SIGNED(-153,11),
TO_SIGNED(-106,11),
TO_SIGNED(-60,11),
TO_SIGNED(-13,11),
TO_SIGNED(34,11),
TO_SIGNED(81,11),
TO_SIGNED(128,11),
TO_SIGNED(174,11),
TO_SIGNED(219,11),
TO_SIGNED(264,11),
TO_SIGNED(307,11),
TO_SIGNED(349,11),
TO_SIGNED(390,11),
TO_SIGNED(430,11),
TO_SIGNED(467,11),
TO_SIGNED(503,11),
TO_SIGNED(537,11),
TO_SIGNED(569,11),
TO_SIGNED(598,11),
TO_SIGNED(625,11),
TO_SIGNED(650,11),
TO_SIGNED(672,11),
TO_SIGNED(692,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(730,11),
TO_SIGNED(718,11),
TO_SIGNED(703,11),
TO_SIGNED(685,11),
TO_SIGNED(665,11),
TO_SIGNED(642,11),
TO_SIGNED(616,11),
TO_SIGNED(588,11),
TO_SIGNED(558,11),
TO_SIGNED(526,11),
TO_SIGNED(491,11),
TO_SIGNED(455,11),
TO_SIGNED(416,11),
TO_SIGNED(376,11),
TO_SIGNED(335,11),
TO_SIGNED(292,11),
TO_SIGNED(248,11),
TO_SIGNED(204,11),
TO_SIGNED(158,11),
TO_SIGNED(112,11),
TO_SIGNED(65,11),
TO_SIGNED(18,11),
TO_SIGNED(-29,11),
TO_SIGNED(-76,11),
TO_SIGNED(-122,11),
TO_SIGNED(-168,11),
TO_SIGNED(-214,11),
TO_SIGNED(-259,11),
TO_SIGNED(-302,11),
TO_SIGNED(-345,11),
TO_SIGNED(-386,11),
TO_SIGNED(-425,11),
TO_SIGNED(-463,11),
TO_SIGNED(-499,11),
TO_SIGNED(-533,11),
TO_SIGNED(-565,11),
TO_SIGNED(-595,11),
TO_SIGNED(-622,11),
TO_SIGNED(-647,11),
TO_SIGNED(-670,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-721,11),
TO_SIGNED(-733,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-720,11),
TO_SIGNED(-705,11),
TO_SIGNED(-688,11),
TO_SIGNED(-667,11),
TO_SIGNED(-645,11),
TO_SIGNED(-619,11),
TO_SIGNED(-592,11),
TO_SIGNED(-562,11),
TO_SIGNED(-529,11),
TO_SIGNED(-495,11),
TO_SIGNED(-459,11),
TO_SIGNED(-421,11),
TO_SIGNED(-381,11),
TO_SIGNED(-340,11),
TO_SIGNED(-297,11),
TO_SIGNED(-254,11),
TO_SIGNED(-209,11),
TO_SIGNED(-163,11),
TO_SIGNED(-117,11),
TO_SIGNED(-70,11),
TO_SIGNED(-24,11),
TO_SIGNED(24,11),
TO_SIGNED(70,11),
TO_SIGNED(117,11),
TO_SIGNED(163,11),
TO_SIGNED(209,11),
TO_SIGNED(254,11),
TO_SIGNED(297,11),
TO_SIGNED(340,11),
TO_SIGNED(381,11),
TO_SIGNED(421,11),
TO_SIGNED(459,11),
TO_SIGNED(495,11),
TO_SIGNED(529,11),
TO_SIGNED(562,11),
TO_SIGNED(592,11),
TO_SIGNED(619,11),
TO_SIGNED(645,11),
TO_SIGNED(667,11),
TO_SIGNED(688,11),
TO_SIGNED(705,11),
TO_SIGNED(720,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(733,11),
TO_SIGNED(721,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(670,11),
TO_SIGNED(647,11),
TO_SIGNED(622,11),
TO_SIGNED(595,11),
TO_SIGNED(565,11),
TO_SIGNED(533,11),
TO_SIGNED(499,11),
TO_SIGNED(463,11),
TO_SIGNED(425,11),
TO_SIGNED(386,11),
TO_SIGNED(345,11),
TO_SIGNED(302,11),
TO_SIGNED(259,11),
TO_SIGNED(214,11),
TO_SIGNED(168,11),
TO_SIGNED(122,11),
TO_SIGNED(76,11),
TO_SIGNED(29,11),
TO_SIGNED(-18,11),
TO_SIGNED(-65,11),
TO_SIGNED(-112,11),
TO_SIGNED(-158,11),
TO_SIGNED(-204,11),
TO_SIGNED(-248,11),
TO_SIGNED(-292,11),
TO_SIGNED(-335,11),
TO_SIGNED(-376,11),
TO_SIGNED(-416,11),
TO_SIGNED(-455,11),
TO_SIGNED(-491,11),
TO_SIGNED(-526,11),
TO_SIGNED(-558,11),
TO_SIGNED(-588,11),
TO_SIGNED(-616,11),
TO_SIGNED(-642,11),
TO_SIGNED(-665,11),
TO_SIGNED(-685,11),
TO_SIGNED(-703,11),
TO_SIGNED(-718,11),
TO_SIGNED(-730,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-692,11),
TO_SIGNED(-672,11),
TO_SIGNED(-650,11),
TO_SIGNED(-625,11),
TO_SIGNED(-598,11),
TO_SIGNED(-569,11),
TO_SIGNED(-537,11),
TO_SIGNED(-503,11),
TO_SIGNED(-467,11),
TO_SIGNED(-430,11),
TO_SIGNED(-390,11),
TO_SIGNED(-349,11),
TO_SIGNED(-307,11),
TO_SIGNED(-264,11),
TO_SIGNED(-219,11),
TO_SIGNED(-174,11),
TO_SIGNED(-128,11),
TO_SIGNED(-81,11),
TO_SIGNED(-34,11),
TO_SIGNED(13,11),
TO_SIGNED(60,11),
TO_SIGNED(106,11),
TO_SIGNED(153,11),
TO_SIGNED(198,11),
TO_SIGNED(243,11),
TO_SIGNED(287,11),
TO_SIGNED(330,11),
TO_SIGNED(372,11),
TO_SIGNED(412,11),
TO_SIGNED(450,11),
TO_SIGNED(487,11),
TO_SIGNED(522,11),
TO_SIGNED(554,11),
TO_SIGNED(585,11),
TO_SIGNED(613,11),
TO_SIGNED(639,11),
TO_SIGNED(662,11),
TO_SIGNED(683,11),
TO_SIGNED(701,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(724,11),
TO_SIGNED(710,11),
TO_SIGNED(694,11),
TO_SIGNED(675,11),
TO_SIGNED(653,11),
TO_SIGNED(628,11),
TO_SIGNED(601,11),
TO_SIGNED(572,11),
TO_SIGNED(541,11),
TO_SIGNED(507,11),
TO_SIGNED(471,11),
TO_SIGNED(434,11),
TO_SIGNED(395,11),
TO_SIGNED(354,11),
TO_SIGNED(312,11),
TO_SIGNED(269,11),
TO_SIGNED(224,11),
TO_SIGNED(179,11),
TO_SIGNED(133,11),
TO_SIGNED(86,11),
TO_SIGNED(40,11),
TO_SIGNED(-7,11),
TO_SIGNED(-54,11),
TO_SIGNED(-101,11),
TO_SIGNED(-148,11),
TO_SIGNED(-193,11),
TO_SIGNED(-238,11),
TO_SIGNED(-282,11),
TO_SIGNED(-325,11),
TO_SIGNED(-367,11),
TO_SIGNED(-407,11),
TO_SIGNED(-446,11),
TO_SIGNED(-483,11),
TO_SIGNED(-518,11),
TO_SIGNED(-551,11),
TO_SIGNED(-582,11),
TO_SIGNED(-610,11),
TO_SIGNED(-636,11),
TO_SIGNED(-660,11),
TO_SIGNED(-681,11),
TO_SIGNED(-699,11),
TO_SIGNED(-715,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-736,11),
TO_SIGNED(-725,11),
TO_SIGNED(-712,11),
TO_SIGNED(-696,11),
TO_SIGNED(-677,11),
TO_SIGNED(-655,11),
TO_SIGNED(-631,11),
TO_SIGNED(-605,11),
TO_SIGNED(-576,11),
TO_SIGNED(-544,11),
TO_SIGNED(-511,11),
TO_SIGNED(-476,11),
TO_SIGNED(-438,11),
TO_SIGNED(-399,11),
TO_SIGNED(-359,11),
TO_SIGNED(-317,11),
TO_SIGNED(-274,11),
TO_SIGNED(-229,11),
TO_SIGNED(-184,11),
TO_SIGNED(-138,11),
TO_SIGNED(-92,11),
TO_SIGNED(-45,11),
TO_SIGNED(2,11),
TO_SIGNED(49,11),
TO_SIGNED(96,11),
TO_SIGNED(142,11),
TO_SIGNED(188,11),
TO_SIGNED(233,11),
TO_SIGNED(277,11),
TO_SIGNED(321,11),
TO_SIGNED(362,11),
TO_SIGNED(403,11),
TO_SIGNED(442,11),
TO_SIGNED(479,11),
TO_SIGNED(514,11),
TO_SIGNED(547,11),
TO_SIGNED(578,11),
TO_SIGNED(607,11),
TO_SIGNED(633,11),
TO_SIGNED(657,11),
TO_SIGNED(679,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(698,11),
TO_SIGNED(679,11),
TO_SIGNED(658,11),
TO_SIGNED(634,11),
TO_SIGNED(608,11),
TO_SIGNED(579,11),
TO_SIGNED(548,11),
TO_SIGNED(515,11),
TO_SIGNED(480,11),
TO_SIGNED(443,11),
TO_SIGNED(404,11),
TO_SIGNED(363,11),
TO_SIGNED(322,11),
TO_SIGNED(278,11),
TO_SIGNED(234,11),
TO_SIGNED(189,11),
TO_SIGNED(143,11),
TO_SIGNED(97,11),
TO_SIGNED(50,11),
TO_SIGNED(3,11),
TO_SIGNED(-44,11),
TO_SIGNED(-91,11),
TO_SIGNED(-137,11),
TO_SIGNED(-183,11),
TO_SIGNED(-228,11),
TO_SIGNED(-273,11),
TO_SIGNED(-316,11),
TO_SIGNED(-358,11),
TO_SIGNED(-398,11),
TO_SIGNED(-437,11),
TO_SIGNED(-475,11),
TO_SIGNED(-510,11),
TO_SIGNED(-544,11),
TO_SIGNED(-575,11),
TO_SIGNED(-604,11),
TO_SIGNED(-631,11),
TO_SIGNED(-655,11),
TO_SIGNED(-676,11),
TO_SIGNED(-695,11),
TO_SIGNED(-712,11),
TO_SIGNED(-725,11),
TO_SIGNED(-736,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-715,11),
TO_SIGNED(-700,11),
TO_SIGNED(-681,11),
TO_SIGNED(-660,11),
TO_SIGNED(-637,11),
TO_SIGNED(-611,11),
TO_SIGNED(-582,11),
TO_SIGNED(-552,11),
TO_SIGNED(-519,11),
TO_SIGNED(-484,11),
TO_SIGNED(-447,11),
TO_SIGNED(-408,11),
TO_SIGNED(-368,11),
TO_SIGNED(-326,11),
TO_SIGNED(-283,11),
TO_SIGNED(-239,11),
TO_SIGNED(-194,11),
TO_SIGNED(-149,11),
TO_SIGNED(-102,11),
TO_SIGNED(-56,11),
TO_SIGNED(-9,11),
TO_SIGNED(38,11),
TO_SIGNED(85,11),
TO_SIGNED(132,11),
TO_SIGNED(178,11),
TO_SIGNED(223,11),
TO_SIGNED(268,11),
TO_SIGNED(311,11),
TO_SIGNED(353,11),
TO_SIGNED(394,11),
TO_SIGNED(433,11),
TO_SIGNED(471,11),
TO_SIGNED(506,11),
TO_SIGNED(540,11),
TO_SIGNED(571,11),
TO_SIGNED(601,11),
TO_SIGNED(628,11),
TO_SIGNED(652,11),
TO_SIGNED(674,11),
TO_SIGNED(693,11),
TO_SIGNED(710,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(739,11),
TO_SIGNED(729,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(684,11),
TO_SIGNED(663,11),
TO_SIGNED(640,11),
TO_SIGNED(614,11),
TO_SIGNED(586,11),
TO_SIGNED(555,11),
TO_SIGNED(523,11),
TO_SIGNED(488,11),
TO_SIGNED(451,11),
TO_SIGNED(413,11),
TO_SIGNED(373,11),
TO_SIGNED(331,11),
TO_SIGNED(288,11),
TO_SIGNED(244,11),
TO_SIGNED(200,11),
TO_SIGNED(154,11),
TO_SIGNED(108,11),
TO_SIGNED(61,11),
TO_SIGNED(14,11),
TO_SIGNED(-33,11),
TO_SIGNED(-80,11),
TO_SIGNED(-127,11),
TO_SIGNED(-173,11),
TO_SIGNED(-218,11),
TO_SIGNED(-263,11),
TO_SIGNED(-306,11),
TO_SIGNED(-348,11),
TO_SIGNED(-389,11),
TO_SIGNED(-429,11),
TO_SIGNED(-466,11),
TO_SIGNED(-502,11),
TO_SIGNED(-536,11),
TO_SIGNED(-568,11),
TO_SIGNED(-598,11),
TO_SIGNED(-625,11),
TO_SIGNED(-650,11),
TO_SIGNED(-672,11),
TO_SIGNED(-691,11),
TO_SIGNED(-708,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-686,11),
TO_SIGNED(-665,11),
TO_SIGNED(-642,11),
TO_SIGNED(-617,11),
TO_SIGNED(-589,11),
TO_SIGNED(-559,11),
TO_SIGNED(-526,11),
TO_SIGNED(-492,11),
TO_SIGNED(-455,11),
TO_SIGNED(-417,11),
TO_SIGNED(-377,11),
TO_SIGNED(-336,11),
TO_SIGNED(-293,11),
TO_SIGNED(-249,11),
TO_SIGNED(-205,11),
TO_SIGNED(-159,11),
TO_SIGNED(-113,11),
TO_SIGNED(-66,11),
TO_SIGNED(-19,11),
TO_SIGNED(28,11),
TO_SIGNED(75,11),
TO_SIGNED(121,11),
TO_SIGNED(167,11),
TO_SIGNED(213,11),
TO_SIGNED(258,11),
TO_SIGNED(301,11),
TO_SIGNED(344,11),
TO_SIGNED(385,11),
TO_SIGNED(424,11),
TO_SIGNED(462,11),
TO_SIGNED(498,11),
TO_SIGNED(532,11),
TO_SIGNED(564,11),
TO_SIGNED(594,11),
TO_SIGNED(622,11),
TO_SIGNED(647,11),
TO_SIGNED(669,11),
TO_SIGNED(689,11),
TO_SIGNED(706,11),
TO_SIGNED(721,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(720,11),
TO_SIGNED(705,11),
TO_SIGNED(688,11),
TO_SIGNED(668,11),
TO_SIGNED(645,11),
TO_SIGNED(620,11),
TO_SIGNED(592,11),
TO_SIGNED(562,11),
TO_SIGNED(530,11),
TO_SIGNED(496,11),
TO_SIGNED(460,11),
TO_SIGNED(422,11),
TO_SIGNED(382,11),
TO_SIGNED(341,11),
TO_SIGNED(298,11),
TO_SIGNED(255,11),
TO_SIGNED(210,11),
TO_SIGNED(164,11),
TO_SIGNED(118,11),
TO_SIGNED(71,11),
TO_SIGNED(25,11),
TO_SIGNED(-22,11),
TO_SIGNED(-69,11),
TO_SIGNED(-116,11),
TO_SIGNED(-162,11),
TO_SIGNED(-208,11),
TO_SIGNED(-252,11),
TO_SIGNED(-296,11),
TO_SIGNED(-339,11),
TO_SIGNED(-380,11),
TO_SIGNED(-420,11),
TO_SIGNED(-458,11),
TO_SIGNED(-494,11),
TO_SIGNED(-529,11),
TO_SIGNED(-561,11),
TO_SIGNED(-591,11),
TO_SIGNED(-619,11),
TO_SIGNED(-644,11),
TO_SIGNED(-667,11),
TO_SIGNED(-687,11),
TO_SIGNED(-705,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-733,11),
TO_SIGNED(-721,11),
TO_SIGNED(-707,11),
TO_SIGNED(-690,11),
TO_SIGNED(-670,11),
TO_SIGNED(-648,11),
TO_SIGNED(-623,11),
TO_SIGNED(-596,11),
TO_SIGNED(-566,11),
TO_SIGNED(-534,11),
TO_SIGNED(-500,11),
TO_SIGNED(-464,11),
TO_SIGNED(-426,11),
TO_SIGNED(-387,11),
TO_SIGNED(-345,11),
TO_SIGNED(-303,11),
TO_SIGNED(-260,11),
TO_SIGNED(-215,11),
TO_SIGNED(-169,11),
TO_SIGNED(-123,11),
TO_SIGNED(-77,11),
TO_SIGNED(-30,11),
TO_SIGNED(17,11),
TO_SIGNED(64,11),
TO_SIGNED(111,11),
TO_SIGNED(157,11),
TO_SIGNED(203,11),
TO_SIGNED(247,11),
TO_SIGNED(291,11),
TO_SIGNED(334,11),
TO_SIGNED(375,11),
TO_SIGNED(415,11),
TO_SIGNED(454,11),
TO_SIGNED(490,11),
TO_SIGNED(525,11),
TO_SIGNED(557,11),
TO_SIGNED(588,11),
TO_SIGNED(616,11),
TO_SIGNED(641,11),
TO_SIGNED(664,11),
TO_SIGNED(685,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(709,11),
TO_SIGNED(692,11),
TO_SIGNED(673,11),
TO_SIGNED(651,11),
TO_SIGNED(626,11),
TO_SIGNED(599,11),
TO_SIGNED(569,11),
TO_SIGNED(538,11),
TO_SIGNED(504,11),
TO_SIGNED(468,11),
TO_SIGNED(430,11),
TO_SIGNED(391,11),
TO_SIGNED(350,11),
TO_SIGNED(308,11),
TO_SIGNED(265,11),
TO_SIGNED(220,11),
TO_SIGNED(175,11),
TO_SIGNED(129,11),
TO_SIGNED(82,11),
TO_SIGNED(35,11),
TO_SIGNED(-12,11),
TO_SIGNED(-59,11),
TO_SIGNED(-105,11),
TO_SIGNED(-152,11),
TO_SIGNED(-197,11),
TO_SIGNED(-242,11),
TO_SIGNED(-286,11),
TO_SIGNED(-329,11),
TO_SIGNED(-371,11),
TO_SIGNED(-411,11),
TO_SIGNED(-449,11),
TO_SIGNED(-486,11),
TO_SIGNED(-521,11),
TO_SIGNED(-554,11),
TO_SIGNED(-584,11),
TO_SIGNED(-613,11),
TO_SIGNED(-639,11),
TO_SIGNED(-662,11),
TO_SIGNED(-683,11),
TO_SIGNED(-701,11),
TO_SIGNED(-716,11),
TO_SIGNED(-729,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-711,11),
TO_SIGNED(-694,11),
TO_SIGNED(-675,11),
TO_SIGNED(-653,11),
TO_SIGNED(-629,11),
TO_SIGNED(-602,11),
TO_SIGNED(-573,11),
TO_SIGNED(-541,11),
TO_SIGNED(-508,11),
TO_SIGNED(-472,11),
TO_SIGNED(-435,11),
TO_SIGNED(-396,11),
TO_SIGNED(-355,11),
TO_SIGNED(-313,11),
TO_SIGNED(-270,11),
TO_SIGNED(-225,11),
TO_SIGNED(-180,11),
TO_SIGNED(-134,11),
TO_SIGNED(-87,11),
TO_SIGNED(-41,11),
TO_SIGNED(6,11),
TO_SIGNED(53,11),
TO_SIGNED(100,11),
TO_SIGNED(147,11),
TO_SIGNED(192,11),
TO_SIGNED(237,11),
TO_SIGNED(281,11),
TO_SIGNED(324,11),
TO_SIGNED(366,11),
TO_SIGNED(406,11),
TO_SIGNED(445,11),
TO_SIGNED(482,11),
TO_SIGNED(517,11),
TO_SIGNED(550,11),
TO_SIGNED(581,11),
TO_SIGNED(610,11),
TO_SIGNED(636,11),
TO_SIGNED(659,11),
TO_SIGNED(681,11),
TO_SIGNED(699,11),
TO_SIGNED(715,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(712,11),
TO_SIGNED(696,11),
TO_SIGNED(677,11),
TO_SIGNED(656,11),
TO_SIGNED(632,11),
TO_SIGNED(605,11),
TO_SIGNED(576,11),
TO_SIGNED(545,11),
TO_SIGNED(512,11),
TO_SIGNED(476,11),
TO_SIGNED(439,11),
TO_SIGNED(400,11),
TO_SIGNED(360,11),
TO_SIGNED(318,11),
TO_SIGNED(275,11),
TO_SIGNED(230,11),
TO_SIGNED(185,11),
TO_SIGNED(139,11),
TO_SIGNED(93,11),
TO_SIGNED(46,11),
TO_SIGNED(-1,11),
TO_SIGNED(-48,11),
TO_SIGNED(-95,11),
TO_SIGNED(-141,11),
TO_SIGNED(-187,11),
TO_SIGNED(-232,11),
TO_SIGNED(-276,11),
TO_SIGNED(-320,11),
TO_SIGNED(-362,11),
TO_SIGNED(-402,11),
TO_SIGNED(-441,11),
TO_SIGNED(-478,11),
TO_SIGNED(-513,11),
TO_SIGNED(-547,11),
TO_SIGNED(-578,11),
TO_SIGNED(-606,11),
TO_SIGNED(-633,11),
TO_SIGNED(-657,11),
TO_SIGNED(-678,11),
TO_SIGNED(-697,11),
TO_SIGNED(-713,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-714,11),
TO_SIGNED(-698,11),
TO_SIGNED(-680,11),
TO_SIGNED(-658,11),
TO_SIGNED(-635,11),
TO_SIGNED(-608,11),
TO_SIGNED(-580,11),
TO_SIGNED(-549,11),
TO_SIGNED(-516,11),
TO_SIGNED(-480,11),
TO_SIGNED(-443,11),
TO_SIGNED(-405,11),
TO_SIGNED(-364,11),
TO_SIGNED(-323,11),
TO_SIGNED(-279,11),
TO_SIGNED(-235,11),
TO_SIGNED(-190,11),
TO_SIGNED(-144,11),
TO_SIGNED(-98,11),
TO_SIGNED(-51,11),
TO_SIGNED(-4,11),
TO_SIGNED(43,11),
TO_SIGNED(90,11),
TO_SIGNED(136,11),
TO_SIGNED(182,11),
TO_SIGNED(227,11),
TO_SIGNED(272,11),
TO_SIGNED(315,11),
TO_SIGNED(357,11),
TO_SIGNED(397,11),
TO_SIGNED(437,11),
TO_SIGNED(474,11),
TO_SIGNED(509,11),
TO_SIGNED(543,11),
TO_SIGNED(574,11),
TO_SIGNED(603,11),
TO_SIGNED(630,11),
TO_SIGNED(654,11),
TO_SIGNED(676,11),
TO_SIGNED(695,11),
TO_SIGNED(711,11),
TO_SIGNED(725,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(716,11),
TO_SIGNED(700,11),
TO_SIGNED(682,11),
TO_SIGNED(661,11),
TO_SIGNED(637,11),
TO_SIGNED(611,11),
TO_SIGNED(583,11),
TO_SIGNED(552,11),
TO_SIGNED(519,11),
TO_SIGNED(485,11),
TO_SIGNED(448,11),
TO_SIGNED(409,11),
TO_SIGNED(369,11),
TO_SIGNED(327,11),
TO_SIGNED(284,11),
TO_SIGNED(240,11),
TO_SIGNED(195,11),
TO_SIGNED(150,11),
TO_SIGNED(103,11),
TO_SIGNED(57,11),
TO_SIGNED(10,11),
TO_SIGNED(-37,11),
TO_SIGNED(-84,11),
TO_SIGNED(-131,11),
TO_SIGNED(-177,11),
TO_SIGNED(-222,11),
TO_SIGNED(-267,11),
TO_SIGNED(-310,11),
TO_SIGNED(-352,11),
TO_SIGNED(-393,11),
TO_SIGNED(-432,11),
TO_SIGNED(-470,11),
TO_SIGNED(-505,11),
TO_SIGNED(-539,11),
TO_SIGNED(-571,11),
TO_SIGNED(-600,11),
TO_SIGNED(-627,11),
TO_SIGNED(-652,11),
TO_SIGNED(-674,11),
TO_SIGNED(-693,11),
TO_SIGNED(-710,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-702,11),
TO_SIGNED(-684,11),
TO_SIGNED(-663,11),
TO_SIGNED(-640,11),
TO_SIGNED(-615,11),
TO_SIGNED(-586,11),
TO_SIGNED(-556,11),
TO_SIGNED(-523,11),
TO_SIGNED(-489,11),
TO_SIGNED(-452,11),
TO_SIGNED(-414,11),
TO_SIGNED(-374,11),
TO_SIGNED(-332,11),
TO_SIGNED(-289,11),
TO_SIGNED(-245,11),
TO_SIGNED(-201,11),
TO_SIGNED(-155,11),
TO_SIGNED(-109,11),
TO_SIGNED(-62,11),
TO_SIGNED(-15,11),
TO_SIGNED(32,11),
TO_SIGNED(79,11),
TO_SIGNED(125,11),
TO_SIGNED(172,11),
TO_SIGNED(217,11),
TO_SIGNED(262,11),
TO_SIGNED(305,11),
TO_SIGNED(347,11),
TO_SIGNED(388,11),
TO_SIGNED(428,11),
TO_SIGNED(466,11),
TO_SIGNED(501,11),
TO_SIGNED(535,11),
TO_SIGNED(567,11),
TO_SIGNED(597,11),
TO_SIGNED(624,11),
TO_SIGNED(649,11),
TO_SIGNED(671,11),
TO_SIGNED(691,11),
TO_SIGNED(708,11),
TO_SIGNED(722,11),
TO_SIGNED(733,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(704,11),
TO_SIGNED(686,11),
TO_SIGNED(666,11),
TO_SIGNED(643,11),
TO_SIGNED(618,11),
TO_SIGNED(590,11),
TO_SIGNED(559,11),
TO_SIGNED(527,11),
TO_SIGNED(493,11),
TO_SIGNED(456,11),
TO_SIGNED(418,11),
TO_SIGNED(378,11),
TO_SIGNED(337,11),
TO_SIGNED(294,11),
TO_SIGNED(250,11),
TO_SIGNED(206,11),
TO_SIGNED(160,11),
TO_SIGNED(114,11),
TO_SIGNED(67,11),
TO_SIGNED(20,11),
TO_SIGNED(-27,11),
TO_SIGNED(-74,11),
TO_SIGNED(-120,11),
TO_SIGNED(-166,11),
TO_SIGNED(-212,11),
TO_SIGNED(-257,11),
TO_SIGNED(-300,11),
TO_SIGNED(-343,11),
TO_SIGNED(-384,11),
TO_SIGNED(-423,11),
TO_SIGNED(-461,11),
TO_SIGNED(-497,11),
TO_SIGNED(-532,11),
TO_SIGNED(-564,11),
TO_SIGNED(-594,11),
TO_SIGNED(-621,11),
TO_SIGNED(-646,11),
TO_SIGNED(-669,11),
TO_SIGNED(-689,11),
TO_SIGNED(-706,11),
TO_SIGNED(-721,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-720,11),
TO_SIGNED(-706,11),
TO_SIGNED(-688,11),
TO_SIGNED(-668,11),
TO_SIGNED(-646,11),
TO_SIGNED(-621,11),
TO_SIGNED(-593,11),
TO_SIGNED(-563,11),
TO_SIGNED(-531,11),
TO_SIGNED(-497,11),
TO_SIGNED(-460,11),
TO_SIGNED(-422,11),
TO_SIGNED(-383,11),
TO_SIGNED(-342,11),
TO_SIGNED(-299,11),
TO_SIGNED(-256,11),
TO_SIGNED(-211,11),
TO_SIGNED(-165,11),
TO_SIGNED(-119,11),
TO_SIGNED(-73,11),
TO_SIGNED(-26,11),
TO_SIGNED(21,11),
TO_SIGNED(68,11),
TO_SIGNED(115,11),
TO_SIGNED(161,11),
TO_SIGNED(207,11),
TO_SIGNED(251,11),
TO_SIGNED(295,11),
TO_SIGNED(338,11),
TO_SIGNED(379,11),
TO_SIGNED(419,11),
TO_SIGNED(457,11),
TO_SIGNED(493,11),
TO_SIGNED(528,11),
TO_SIGNED(560,11),
TO_SIGNED(590,11),
TO_SIGNED(618,11),
TO_SIGNED(644,11),
TO_SIGNED(666,11),
TO_SIGNED(687,11),
TO_SIGNED(704,11),
TO_SIGNED(719,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(671,11),
TO_SIGNED(648,11),
TO_SIGNED(624,11),
TO_SIGNED(596,11),
TO_SIGNED(567,11),
TO_SIGNED(535,11),
TO_SIGNED(501,11),
TO_SIGNED(465,11),
TO_SIGNED(427,11),
TO_SIGNED(387,11),
TO_SIGNED(346,11),
TO_SIGNED(304,11),
TO_SIGNED(261,11),
TO_SIGNED(216,11),
TO_SIGNED(171,11),
TO_SIGNED(124,11),
TO_SIGNED(78,11),
TO_SIGNED(31,11),
TO_SIGNED(-16,11),
TO_SIGNED(-63,11),
TO_SIGNED(-110,11),
TO_SIGNED(-156,11),
TO_SIGNED(-202,11),
TO_SIGNED(-246,11),
TO_SIGNED(-290,11),
TO_SIGNED(-333,11),
TO_SIGNED(-375,11),
TO_SIGNED(-415,11),
TO_SIGNED(-453,11),
TO_SIGNED(-489,11),
TO_SIGNED(-524,11),
TO_SIGNED(-557,11),
TO_SIGNED(-587,11),
TO_SIGNED(-615,11),
TO_SIGNED(-641,11),
TO_SIGNED(-664,11),
TO_SIGNED(-685,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-730,11),
TO_SIGNED(-739,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-693,11),
TO_SIGNED(-673,11),
TO_SIGNED(-651,11),
TO_SIGNED(-627,11),
TO_SIGNED(-599,11),
TO_SIGNED(-570,11),
TO_SIGNED(-538,11),
TO_SIGNED(-505,11),
TO_SIGNED(-469,11),
TO_SIGNED(-431,11),
TO_SIGNED(-392,11),
TO_SIGNED(-351,11),
TO_SIGNED(-309,11),
TO_SIGNED(-266,11),
TO_SIGNED(-221,11),
TO_SIGNED(-176,11),
TO_SIGNED(-130,11),
TO_SIGNED(-83,11),
TO_SIGNED(-36,11),
TO_SIGNED(11,11),
TO_SIGNED(58,11),
TO_SIGNED(104,11),
TO_SIGNED(151,11),
TO_SIGNED(196,11),
TO_SIGNED(241,11),
TO_SIGNED(285,11),
TO_SIGNED(328,11),
TO_SIGNED(370,11),
TO_SIGNED(410,11),
TO_SIGNED(449,11),
TO_SIGNED(485,11),
TO_SIGNED(520,11),
TO_SIGNED(553,11),
TO_SIGNED(584,11),
TO_SIGNED(612,11),
TO_SIGNED(638,11),
TO_SIGNED(661,11),
TO_SIGNED(682,11),
TO_SIGNED(700,11),
TO_SIGNED(716,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(725,11),
TO_SIGNED(711,11),
TO_SIGNED(695,11),
TO_SIGNED(675,11),
TO_SIGNED(654,11),
TO_SIGNED(629,11),
TO_SIGNED(603,11),
TO_SIGNED(574,11),
TO_SIGNED(542,11),
TO_SIGNED(509,11),
TO_SIGNED(473,11),
TO_SIGNED(436,11),
TO_SIGNED(397,11),
TO_SIGNED(356,11),
TO_SIGNED(314,11),
TO_SIGNED(271,11),
TO_SIGNED(226,11),
TO_SIGNED(181,11),
TO_SIGNED(135,11),
TO_SIGNED(88,11),
TO_SIGNED(42,11),
TO_SIGNED(-5,11),
TO_SIGNED(-52,11),
TO_SIGNED(-99,11),
TO_SIGNED(-145,11),
TO_SIGNED(-191,11),
TO_SIGNED(-236,11),
TO_SIGNED(-280,11),
TO_SIGNED(-323,11),
TO_SIGNED(-365,11),
TO_SIGNED(-406,11),
TO_SIGNED(-444,11),
TO_SIGNED(-481,11),
TO_SIGNED(-516,11),
TO_SIGNED(-549,11),
TO_SIGNED(-580,11),
TO_SIGNED(-609,11),
TO_SIGNED(-635,11),
TO_SIGNED(-659,11),
TO_SIGNED(-680,11),
TO_SIGNED(-699,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-736,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-678,11),
TO_SIGNED(-656,11),
TO_SIGNED(-632,11),
TO_SIGNED(-606,11),
TO_SIGNED(-577,11),
TO_SIGNED(-546,11),
TO_SIGNED(-512,11),
TO_SIGNED(-477,11),
TO_SIGNED(-440,11),
TO_SIGNED(-401,11),
TO_SIGNED(-361,11),
TO_SIGNED(-319,11),
TO_SIGNED(-275,11),
TO_SIGNED(-231,11),
TO_SIGNED(-186,11),
TO_SIGNED(-140,11),
TO_SIGNED(-94,11),
TO_SIGNED(-47,11),
TO_SIGNED(0,11),
TO_SIGNED(47,11),
TO_SIGNED(94,11),
TO_SIGNED(140,11),
TO_SIGNED(186,11),
TO_SIGNED(231,11),
TO_SIGNED(275,11),
TO_SIGNED(319,11),
TO_SIGNED(361,11),
TO_SIGNED(401,11),
TO_SIGNED(440,11),
TO_SIGNED(477,11),
TO_SIGNED(512,11),
TO_SIGNED(546,11),
TO_SIGNED(577,11),
TO_SIGNED(606,11),
TO_SIGNED(632,11),
TO_SIGNED(656,11),
TO_SIGNED(678,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(736,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(699,11),
TO_SIGNED(680,11),
TO_SIGNED(659,11),
TO_SIGNED(635,11),
TO_SIGNED(609,11),
TO_SIGNED(580,11),
TO_SIGNED(549,11),
TO_SIGNED(516,11),
TO_SIGNED(481,11),
TO_SIGNED(444,11),
TO_SIGNED(406,11),
TO_SIGNED(365,11),
TO_SIGNED(323,11),
TO_SIGNED(280,11),
TO_SIGNED(236,11),
TO_SIGNED(191,11),
TO_SIGNED(145,11),
TO_SIGNED(99,11),
TO_SIGNED(52,11),
TO_SIGNED(5,11),
TO_SIGNED(-42,11),
TO_SIGNED(-88,11),
TO_SIGNED(-135,11),
TO_SIGNED(-181,11),
TO_SIGNED(-226,11),
TO_SIGNED(-271,11),
TO_SIGNED(-314,11),
TO_SIGNED(-356,11),
TO_SIGNED(-397,11),
TO_SIGNED(-436,11),
TO_SIGNED(-473,11),
TO_SIGNED(-509,11),
TO_SIGNED(-542,11),
TO_SIGNED(-574,11),
TO_SIGNED(-603,11),
TO_SIGNED(-629,11),
TO_SIGNED(-654,11),
TO_SIGNED(-675,11),
TO_SIGNED(-695,11),
TO_SIGNED(-711,11),
TO_SIGNED(-725,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-716,11),
TO_SIGNED(-700,11),
TO_SIGNED(-682,11),
TO_SIGNED(-661,11),
TO_SIGNED(-638,11),
TO_SIGNED(-612,11),
TO_SIGNED(-584,11),
TO_SIGNED(-553,11),
TO_SIGNED(-520,11),
TO_SIGNED(-485,11),
TO_SIGNED(-449,11),
TO_SIGNED(-410,11),
TO_SIGNED(-370,11),
TO_SIGNED(-328,11),
TO_SIGNED(-285,11),
TO_SIGNED(-241,11),
TO_SIGNED(-196,11),
TO_SIGNED(-151,11),
TO_SIGNED(-104,11),
TO_SIGNED(-58,11),
TO_SIGNED(-11,11),
TO_SIGNED(36,11),
TO_SIGNED(83,11),
TO_SIGNED(130,11),
TO_SIGNED(176,11),
TO_SIGNED(221,11),
TO_SIGNED(266,11),
TO_SIGNED(309,11),
TO_SIGNED(351,11),
TO_SIGNED(392,11),
TO_SIGNED(431,11),
TO_SIGNED(469,11),
TO_SIGNED(505,11),
TO_SIGNED(538,11),
TO_SIGNED(570,11),
TO_SIGNED(599,11),
TO_SIGNED(627,11),
TO_SIGNED(651,11),
TO_SIGNED(673,11),
TO_SIGNED(693,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(739,11),
TO_SIGNED(730,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(685,11),
TO_SIGNED(664,11),
TO_SIGNED(641,11),
TO_SIGNED(615,11),
TO_SIGNED(587,11),
TO_SIGNED(557,11),
TO_SIGNED(524,11),
TO_SIGNED(489,11),
TO_SIGNED(453,11),
TO_SIGNED(415,11),
TO_SIGNED(375,11),
TO_SIGNED(333,11),
TO_SIGNED(290,11),
TO_SIGNED(246,11),
TO_SIGNED(202,11),
TO_SIGNED(156,11),
TO_SIGNED(110,11),
TO_SIGNED(63,11),
TO_SIGNED(16,11),
TO_SIGNED(-31,11),
TO_SIGNED(-78,11),
TO_SIGNED(-124,11),
TO_SIGNED(-171,11),
TO_SIGNED(-216,11),
TO_SIGNED(-261,11),
TO_SIGNED(-304,11),
TO_SIGNED(-346,11),
TO_SIGNED(-387,11),
TO_SIGNED(-427,11),
TO_SIGNED(-465,11),
TO_SIGNED(-501,11),
TO_SIGNED(-535,11),
TO_SIGNED(-567,11),
TO_SIGNED(-596,11),
TO_SIGNED(-624,11),
TO_SIGNED(-648,11),
TO_SIGNED(-671,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-719,11),
TO_SIGNED(-704,11),
TO_SIGNED(-687,11),
TO_SIGNED(-666,11),
TO_SIGNED(-644,11),
TO_SIGNED(-618,11),
TO_SIGNED(-590,11),
TO_SIGNED(-560,11),
TO_SIGNED(-528,11),
TO_SIGNED(-493,11),
TO_SIGNED(-457,11),
TO_SIGNED(-419,11),
TO_SIGNED(-379,11),
TO_SIGNED(-338,11),
TO_SIGNED(-295,11),
TO_SIGNED(-251,11),
TO_SIGNED(-207,11),
TO_SIGNED(-161,11),
TO_SIGNED(-115,11),
TO_SIGNED(-68,11),
TO_SIGNED(-21,11),
TO_SIGNED(26,11),
TO_SIGNED(73,11),
TO_SIGNED(119,11),
TO_SIGNED(165,11),
TO_SIGNED(211,11),
TO_SIGNED(256,11),
TO_SIGNED(299,11),
TO_SIGNED(342,11),
TO_SIGNED(383,11),
TO_SIGNED(422,11),
TO_SIGNED(460,11),
TO_SIGNED(497,11),
TO_SIGNED(531,11),
TO_SIGNED(563,11),
TO_SIGNED(593,11),
TO_SIGNED(621,11),
TO_SIGNED(646,11),
TO_SIGNED(668,11),
TO_SIGNED(688,11),
TO_SIGNED(706,11),
TO_SIGNED(720,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(721,11),
TO_SIGNED(706,11),
TO_SIGNED(689,11),
TO_SIGNED(669,11),
TO_SIGNED(646,11),
TO_SIGNED(621,11),
TO_SIGNED(594,11),
TO_SIGNED(564,11),
TO_SIGNED(532,11),
TO_SIGNED(497,11),
TO_SIGNED(461,11),
TO_SIGNED(423,11),
TO_SIGNED(384,11),
TO_SIGNED(343,11),
TO_SIGNED(300,11),
TO_SIGNED(257,11),
TO_SIGNED(212,11),
TO_SIGNED(166,11),
TO_SIGNED(120,11),
TO_SIGNED(74,11),
TO_SIGNED(27,11),
TO_SIGNED(-20,11),
TO_SIGNED(-67,11),
TO_SIGNED(-114,11),
TO_SIGNED(-160,11),
TO_SIGNED(-206,11),
TO_SIGNED(-250,11),
TO_SIGNED(-294,11),
TO_SIGNED(-337,11),
TO_SIGNED(-378,11),
TO_SIGNED(-418,11),
TO_SIGNED(-456,11),
TO_SIGNED(-493,11),
TO_SIGNED(-527,11),
TO_SIGNED(-559,11),
TO_SIGNED(-590,11),
TO_SIGNED(-618,11),
TO_SIGNED(-643,11),
TO_SIGNED(-666,11),
TO_SIGNED(-686,11),
TO_SIGNED(-704,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-733,11),
TO_SIGNED(-722,11),
TO_SIGNED(-708,11),
TO_SIGNED(-691,11),
TO_SIGNED(-671,11),
TO_SIGNED(-649,11),
TO_SIGNED(-624,11),
TO_SIGNED(-597,11),
TO_SIGNED(-567,11),
TO_SIGNED(-535,11),
TO_SIGNED(-501,11),
TO_SIGNED(-466,11),
TO_SIGNED(-428,11),
TO_SIGNED(-388,11),
TO_SIGNED(-347,11),
TO_SIGNED(-305,11),
TO_SIGNED(-262,11),
TO_SIGNED(-217,11),
TO_SIGNED(-172,11),
TO_SIGNED(-125,11),
TO_SIGNED(-79,11),
TO_SIGNED(-32,11),
TO_SIGNED(15,11),
TO_SIGNED(62,11),
TO_SIGNED(109,11),
TO_SIGNED(155,11),
TO_SIGNED(201,11),
TO_SIGNED(245,11),
TO_SIGNED(289,11),
TO_SIGNED(332,11),
TO_SIGNED(374,11),
TO_SIGNED(414,11),
TO_SIGNED(452,11),
TO_SIGNED(489,11),
TO_SIGNED(523,11),
TO_SIGNED(556,11),
TO_SIGNED(586,11),
TO_SIGNED(615,11),
TO_SIGNED(640,11),
TO_SIGNED(663,11),
TO_SIGNED(684,11),
TO_SIGNED(702,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(710,11),
TO_SIGNED(693,11),
TO_SIGNED(674,11),
TO_SIGNED(652,11),
TO_SIGNED(627,11),
TO_SIGNED(600,11),
TO_SIGNED(571,11),
TO_SIGNED(539,11),
TO_SIGNED(505,11),
TO_SIGNED(470,11),
TO_SIGNED(432,11),
TO_SIGNED(393,11),
TO_SIGNED(352,11),
TO_SIGNED(310,11),
TO_SIGNED(267,11),
TO_SIGNED(222,11),
TO_SIGNED(177,11),
TO_SIGNED(131,11),
TO_SIGNED(84,11),
TO_SIGNED(37,11),
TO_SIGNED(-10,11),
TO_SIGNED(-57,11),
TO_SIGNED(-103,11),
TO_SIGNED(-150,11),
TO_SIGNED(-195,11),
TO_SIGNED(-240,11),
TO_SIGNED(-284,11),
TO_SIGNED(-327,11),
TO_SIGNED(-369,11),
TO_SIGNED(-409,11),
TO_SIGNED(-448,11),
TO_SIGNED(-485,11),
TO_SIGNED(-519,11),
TO_SIGNED(-552,11),
TO_SIGNED(-583,11),
TO_SIGNED(-611,11),
TO_SIGNED(-637,11),
TO_SIGNED(-661,11),
TO_SIGNED(-682,11),
TO_SIGNED(-700,11),
TO_SIGNED(-716,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-725,11),
TO_SIGNED(-711,11),
TO_SIGNED(-695,11),
TO_SIGNED(-676,11),
TO_SIGNED(-654,11),
TO_SIGNED(-630,11),
TO_SIGNED(-603,11),
TO_SIGNED(-574,11),
TO_SIGNED(-543,11),
TO_SIGNED(-509,11),
TO_SIGNED(-474,11),
TO_SIGNED(-437,11),
TO_SIGNED(-397,11),
TO_SIGNED(-357,11),
TO_SIGNED(-315,11),
TO_SIGNED(-272,11),
TO_SIGNED(-227,11),
TO_SIGNED(-182,11),
TO_SIGNED(-136,11),
TO_SIGNED(-90,11),
TO_SIGNED(-43,11),
TO_SIGNED(4,11),
TO_SIGNED(51,11),
TO_SIGNED(98,11),
TO_SIGNED(144,11),
TO_SIGNED(190,11),
TO_SIGNED(235,11),
TO_SIGNED(279,11),
TO_SIGNED(323,11),
TO_SIGNED(364,11),
TO_SIGNED(405,11),
TO_SIGNED(443,11),
TO_SIGNED(480,11),
TO_SIGNED(516,11),
TO_SIGNED(549,11),
TO_SIGNED(580,11),
TO_SIGNED(608,11),
TO_SIGNED(635,11),
TO_SIGNED(658,11),
TO_SIGNED(680,11),
TO_SIGNED(698,11),
TO_SIGNED(714,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(713,11),
TO_SIGNED(697,11),
TO_SIGNED(678,11),
TO_SIGNED(657,11),
TO_SIGNED(633,11),
TO_SIGNED(606,11),
TO_SIGNED(578,11),
TO_SIGNED(547,11),
TO_SIGNED(513,11),
TO_SIGNED(478,11),
TO_SIGNED(441,11),
TO_SIGNED(402,11),
TO_SIGNED(362,11),
TO_SIGNED(320,11),
TO_SIGNED(276,11),
TO_SIGNED(232,11),
TO_SIGNED(187,11),
TO_SIGNED(141,11),
TO_SIGNED(95,11),
TO_SIGNED(48,11),
TO_SIGNED(1,11),
TO_SIGNED(-46,11),
TO_SIGNED(-93,11),
TO_SIGNED(-139,11),
TO_SIGNED(-185,11),
TO_SIGNED(-230,11),
TO_SIGNED(-275,11),
TO_SIGNED(-318,11),
TO_SIGNED(-360,11),
TO_SIGNED(-400,11),
TO_SIGNED(-439,11),
TO_SIGNED(-476,11),
TO_SIGNED(-512,11),
TO_SIGNED(-545,11),
TO_SIGNED(-576,11),
TO_SIGNED(-605,11),
TO_SIGNED(-632,11),
TO_SIGNED(-656,11),
TO_SIGNED(-677,11),
TO_SIGNED(-696,11),
TO_SIGNED(-712,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-715,11),
TO_SIGNED(-699,11),
TO_SIGNED(-681,11),
TO_SIGNED(-659,11),
TO_SIGNED(-636,11),
TO_SIGNED(-610,11),
TO_SIGNED(-581,11),
TO_SIGNED(-550,11),
TO_SIGNED(-517,11),
TO_SIGNED(-482,11),
TO_SIGNED(-445,11),
TO_SIGNED(-406,11),
TO_SIGNED(-366,11),
TO_SIGNED(-324,11),
TO_SIGNED(-281,11),
TO_SIGNED(-237,11),
TO_SIGNED(-192,11),
TO_SIGNED(-147,11),
TO_SIGNED(-100,11),
TO_SIGNED(-53,11),
TO_SIGNED(-6,11),
TO_SIGNED(41,11),
TO_SIGNED(87,11),
TO_SIGNED(134,11),
TO_SIGNED(180,11),
TO_SIGNED(225,11),
TO_SIGNED(270,11),
TO_SIGNED(313,11),
TO_SIGNED(355,11),
TO_SIGNED(396,11),
TO_SIGNED(435,11),
TO_SIGNED(472,11),
TO_SIGNED(508,11),
TO_SIGNED(541,11),
TO_SIGNED(573,11),
TO_SIGNED(602,11),
TO_SIGNED(629,11),
TO_SIGNED(653,11),
TO_SIGNED(675,11),
TO_SIGNED(694,11),
TO_SIGNED(711,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(729,11),
TO_SIGNED(716,11),
TO_SIGNED(701,11),
TO_SIGNED(683,11),
TO_SIGNED(662,11),
TO_SIGNED(639,11),
TO_SIGNED(613,11),
TO_SIGNED(584,11),
TO_SIGNED(554,11),
TO_SIGNED(521,11),
TO_SIGNED(486,11),
TO_SIGNED(449,11),
TO_SIGNED(411,11),
TO_SIGNED(371,11),
TO_SIGNED(329,11),
TO_SIGNED(286,11),
TO_SIGNED(242,11),
TO_SIGNED(197,11),
TO_SIGNED(152,11),
TO_SIGNED(105,11),
TO_SIGNED(59,11),
TO_SIGNED(12,11),
TO_SIGNED(-35,11),
TO_SIGNED(-82,11),
TO_SIGNED(-129,11),
TO_SIGNED(-175,11),
TO_SIGNED(-220,11),
TO_SIGNED(-265,11),
TO_SIGNED(-308,11),
TO_SIGNED(-350,11),
TO_SIGNED(-391,11),
TO_SIGNED(-430,11),
TO_SIGNED(-468,11),
TO_SIGNED(-504,11),
TO_SIGNED(-538,11),
TO_SIGNED(-569,11),
TO_SIGNED(-599,11),
TO_SIGNED(-626,11),
TO_SIGNED(-651,11),
TO_SIGNED(-673,11),
TO_SIGNED(-692,11),
TO_SIGNED(-709,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-685,11),
TO_SIGNED(-664,11),
TO_SIGNED(-641,11),
TO_SIGNED(-616,11),
TO_SIGNED(-588,11),
TO_SIGNED(-557,11),
TO_SIGNED(-525,11),
TO_SIGNED(-490,11),
TO_SIGNED(-454,11),
TO_SIGNED(-415,11),
TO_SIGNED(-375,11),
TO_SIGNED(-334,11),
TO_SIGNED(-291,11),
TO_SIGNED(-247,11),
TO_SIGNED(-203,11),
TO_SIGNED(-157,11),
TO_SIGNED(-111,11),
TO_SIGNED(-64,11),
TO_SIGNED(-17,11),
TO_SIGNED(30,11),
TO_SIGNED(77,11),
TO_SIGNED(123,11),
TO_SIGNED(169,11),
TO_SIGNED(215,11),
TO_SIGNED(260,11),
TO_SIGNED(303,11),
TO_SIGNED(345,11),
TO_SIGNED(387,11),
TO_SIGNED(426,11),
TO_SIGNED(464,11),
TO_SIGNED(500,11),
TO_SIGNED(534,11),
TO_SIGNED(566,11),
TO_SIGNED(596,11),
TO_SIGNED(623,11),
TO_SIGNED(648,11),
TO_SIGNED(670,11),
TO_SIGNED(690,11),
TO_SIGNED(707,11),
TO_SIGNED(721,11),
TO_SIGNED(733,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(705,11),
TO_SIGNED(687,11),
TO_SIGNED(667,11),
TO_SIGNED(644,11),
TO_SIGNED(619,11),
TO_SIGNED(591,11),
TO_SIGNED(561,11),
TO_SIGNED(529,11),
TO_SIGNED(494,11),
TO_SIGNED(458,11),
TO_SIGNED(420,11),
TO_SIGNED(380,11),
TO_SIGNED(339,11),
TO_SIGNED(296,11),
TO_SIGNED(252,11),
TO_SIGNED(208,11),
TO_SIGNED(162,11),
TO_SIGNED(116,11),
TO_SIGNED(69,11),
TO_SIGNED(22,11),
TO_SIGNED(-25,11),
TO_SIGNED(-71,11),
TO_SIGNED(-118,11),
TO_SIGNED(-164,11),
TO_SIGNED(-210,11),
TO_SIGNED(-255,11),
TO_SIGNED(-298,11),
TO_SIGNED(-341,11),
TO_SIGNED(-382,11),
TO_SIGNED(-422,11),
TO_SIGNED(-460,11),
TO_SIGNED(-496,11),
TO_SIGNED(-530,11),
TO_SIGNED(-562,11),
TO_SIGNED(-592,11),
TO_SIGNED(-620,11),
TO_SIGNED(-645,11),
TO_SIGNED(-668,11),
TO_SIGNED(-688,11),
TO_SIGNED(-705,11),
TO_SIGNED(-720,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-721,11),
TO_SIGNED(-706,11),
TO_SIGNED(-689,11),
TO_SIGNED(-669,11),
TO_SIGNED(-647,11),
TO_SIGNED(-622,11),
TO_SIGNED(-594,11),
TO_SIGNED(-564,11),
TO_SIGNED(-532,11),
TO_SIGNED(-498,11),
TO_SIGNED(-462,11),
TO_SIGNED(-424,11),
TO_SIGNED(-385,11),
TO_SIGNED(-344,11),
TO_SIGNED(-301,11),
TO_SIGNED(-258,11),
TO_SIGNED(-213,11),
TO_SIGNED(-167,11),
TO_SIGNED(-121,11),
TO_SIGNED(-75,11),
TO_SIGNED(-28,11),
TO_SIGNED(19,11),
TO_SIGNED(66,11),
TO_SIGNED(113,11),
TO_SIGNED(159,11),
TO_SIGNED(205,11),
TO_SIGNED(249,11),
TO_SIGNED(293,11),
TO_SIGNED(336,11),
TO_SIGNED(377,11),
TO_SIGNED(417,11),
TO_SIGNED(455,11),
TO_SIGNED(492,11),
TO_SIGNED(526,11),
TO_SIGNED(559,11),
TO_SIGNED(589,11),
TO_SIGNED(617,11),
TO_SIGNED(642,11),
TO_SIGNED(665,11),
TO_SIGNED(686,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(708,11),
TO_SIGNED(691,11),
TO_SIGNED(672,11),
TO_SIGNED(650,11),
TO_SIGNED(625,11),
TO_SIGNED(598,11),
TO_SIGNED(568,11),
TO_SIGNED(536,11),
TO_SIGNED(502,11),
TO_SIGNED(466,11),
TO_SIGNED(429,11),
TO_SIGNED(389,11),
TO_SIGNED(348,11),
TO_SIGNED(306,11),
TO_SIGNED(263,11),
TO_SIGNED(218,11),
TO_SIGNED(173,11),
TO_SIGNED(127,11),
TO_SIGNED(80,11),
TO_SIGNED(33,11),
TO_SIGNED(-14,11),
TO_SIGNED(-61,11),
TO_SIGNED(-108,11),
TO_SIGNED(-154,11),
TO_SIGNED(-200,11),
TO_SIGNED(-244,11),
TO_SIGNED(-288,11),
TO_SIGNED(-331,11),
TO_SIGNED(-373,11),
TO_SIGNED(-413,11),
TO_SIGNED(-451,11),
TO_SIGNED(-488,11),
TO_SIGNED(-523,11),
TO_SIGNED(-555,11),
TO_SIGNED(-586,11),
TO_SIGNED(-614,11),
TO_SIGNED(-640,11),
TO_SIGNED(-663,11),
TO_SIGNED(-684,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-729,11),
TO_SIGNED(-739,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-710,11),
TO_SIGNED(-693,11),
TO_SIGNED(-674,11),
TO_SIGNED(-652,11),
TO_SIGNED(-628,11),
TO_SIGNED(-601,11),
TO_SIGNED(-571,11),
TO_SIGNED(-540,11),
TO_SIGNED(-506,11),
TO_SIGNED(-471,11),
TO_SIGNED(-433,11),
TO_SIGNED(-394,11),
TO_SIGNED(-353,11),
TO_SIGNED(-311,11),
TO_SIGNED(-268,11),
TO_SIGNED(-223,11),
TO_SIGNED(-178,11),
TO_SIGNED(-132,11),
TO_SIGNED(-85,11),
TO_SIGNED(-38,11),
TO_SIGNED(9,11),
TO_SIGNED(56,11),
TO_SIGNED(102,11),
TO_SIGNED(149,11),
TO_SIGNED(194,11),
TO_SIGNED(239,11),
TO_SIGNED(283,11),
TO_SIGNED(326,11),
TO_SIGNED(368,11),
TO_SIGNED(408,11),
TO_SIGNED(447,11),
TO_SIGNED(484,11),
TO_SIGNED(519,11),
TO_SIGNED(552,11),
TO_SIGNED(582,11),
TO_SIGNED(611,11),
TO_SIGNED(637,11),
TO_SIGNED(660,11),
TO_SIGNED(681,11),
TO_SIGNED(700,11),
TO_SIGNED(715,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(736,11),
TO_SIGNED(725,11),
TO_SIGNED(712,11),
TO_SIGNED(695,11),
TO_SIGNED(676,11),
TO_SIGNED(655,11),
TO_SIGNED(631,11),
TO_SIGNED(604,11),
TO_SIGNED(575,11),
TO_SIGNED(544,11),
TO_SIGNED(510,11),
TO_SIGNED(475,11),
TO_SIGNED(437,11),
TO_SIGNED(398,11),
TO_SIGNED(358,11),
TO_SIGNED(316,11),
TO_SIGNED(273,11),
TO_SIGNED(228,11),
TO_SIGNED(183,11),
TO_SIGNED(137,11),
TO_SIGNED(91,11),
TO_SIGNED(44,11),
TO_SIGNED(-3,11),
TO_SIGNED(-50,11),
TO_SIGNED(-97,11),
TO_SIGNED(-143,11),
TO_SIGNED(-189,11),
TO_SIGNED(-234,11),
TO_SIGNED(-278,11),
TO_SIGNED(-322,11),
TO_SIGNED(-363,11),
TO_SIGNED(-404,11),
TO_SIGNED(-443,11),
TO_SIGNED(-480,11),
TO_SIGNED(-515,11),
TO_SIGNED(-548,11),
TO_SIGNED(-579,11),
TO_SIGNED(-608,11),
TO_SIGNED(-634,11),
TO_SIGNED(-658,11),
TO_SIGNED(-679,11),
TO_SIGNED(-698,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-679,11),
TO_SIGNED(-657,11),
TO_SIGNED(-633,11),
TO_SIGNED(-607,11),
TO_SIGNED(-578,11),
TO_SIGNED(-547,11),
TO_SIGNED(-514,11),
TO_SIGNED(-479,11),
TO_SIGNED(-442,11),
TO_SIGNED(-403,11),
TO_SIGNED(-362,11),
TO_SIGNED(-321,11),
TO_SIGNED(-277,11),
TO_SIGNED(-233,11),
TO_SIGNED(-188,11),
TO_SIGNED(-142,11),
TO_SIGNED(-96,11),
TO_SIGNED(-49,11),
TO_SIGNED(-2,11),
TO_SIGNED(45,11),
TO_SIGNED(92,11),
TO_SIGNED(138,11),
TO_SIGNED(184,11),
TO_SIGNED(229,11),
TO_SIGNED(274,11),
TO_SIGNED(317,11),
TO_SIGNED(359,11),
TO_SIGNED(399,11),
TO_SIGNED(438,11),
TO_SIGNED(476,11),
TO_SIGNED(511,11),
TO_SIGNED(544,11),
TO_SIGNED(576,11),
TO_SIGNED(605,11),
TO_SIGNED(631,11),
TO_SIGNED(655,11),
TO_SIGNED(677,11),
TO_SIGNED(696,11),
TO_SIGNED(712,11),
TO_SIGNED(725,11),
TO_SIGNED(736,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(715,11),
TO_SIGNED(699,11),
TO_SIGNED(681,11),
TO_SIGNED(660,11),
TO_SIGNED(636,11),
TO_SIGNED(610,11),
TO_SIGNED(582,11),
TO_SIGNED(551,11),
TO_SIGNED(518,11),
TO_SIGNED(483,11),
TO_SIGNED(446,11),
TO_SIGNED(407,11),
TO_SIGNED(367,11),
TO_SIGNED(325,11),
TO_SIGNED(282,11),
TO_SIGNED(238,11),
TO_SIGNED(193,11),
TO_SIGNED(148,11),
TO_SIGNED(101,11),
TO_SIGNED(54,11),
TO_SIGNED(7,11),
TO_SIGNED(-40,11),
TO_SIGNED(-86,11),
TO_SIGNED(-133,11),
TO_SIGNED(-179,11),
TO_SIGNED(-224,11),
TO_SIGNED(-269,11),
TO_SIGNED(-312,11),
TO_SIGNED(-354,11),
TO_SIGNED(-395,11),
TO_SIGNED(-434,11),
TO_SIGNED(-471,11),
TO_SIGNED(-507,11),
TO_SIGNED(-541,11),
TO_SIGNED(-572,11),
TO_SIGNED(-601,11),
TO_SIGNED(-628,11),
TO_SIGNED(-653,11),
TO_SIGNED(-675,11),
TO_SIGNED(-694,11),
TO_SIGNED(-710,11),
TO_SIGNED(-724,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-701,11),
TO_SIGNED(-683,11),
TO_SIGNED(-662,11),
TO_SIGNED(-639,11),
TO_SIGNED(-613,11),
TO_SIGNED(-585,11),
TO_SIGNED(-554,11),
TO_SIGNED(-522,11),
TO_SIGNED(-487,11),
TO_SIGNED(-450,11),
TO_SIGNED(-412,11),
TO_SIGNED(-372,11),
TO_SIGNED(-330,11),
TO_SIGNED(-287,11),
TO_SIGNED(-243,11),
TO_SIGNED(-198,11),
TO_SIGNED(-153,11),
TO_SIGNED(-106,11),
TO_SIGNED(-60,11),
TO_SIGNED(-13,11),
TO_SIGNED(34,11),
TO_SIGNED(81,11),
TO_SIGNED(128,11),
TO_SIGNED(174,11),
TO_SIGNED(219,11),
TO_SIGNED(264,11),
TO_SIGNED(307,11),
TO_SIGNED(349,11),
TO_SIGNED(390,11),
TO_SIGNED(430,11),
TO_SIGNED(467,11),
TO_SIGNED(503,11),
TO_SIGNED(537,11),
TO_SIGNED(569,11),
TO_SIGNED(598,11),
TO_SIGNED(625,11),
TO_SIGNED(650,11),
TO_SIGNED(672,11),
TO_SIGNED(692,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(730,11),
TO_SIGNED(718,11),
TO_SIGNED(703,11),
TO_SIGNED(685,11),
TO_SIGNED(665,11),
TO_SIGNED(642,11),
TO_SIGNED(616,11),
TO_SIGNED(588,11),
TO_SIGNED(558,11),
TO_SIGNED(526,11),
TO_SIGNED(491,11),
TO_SIGNED(455,11),
TO_SIGNED(416,11),
TO_SIGNED(376,11),
TO_SIGNED(335,11),
TO_SIGNED(292,11),
TO_SIGNED(248,11),
TO_SIGNED(204,11),
TO_SIGNED(158,11),
TO_SIGNED(112,11),
TO_SIGNED(65,11),
TO_SIGNED(18,11),
TO_SIGNED(-29,11),
TO_SIGNED(-76,11),
TO_SIGNED(-122,11),
TO_SIGNED(-168,11),
TO_SIGNED(-214,11),
TO_SIGNED(-259,11),
TO_SIGNED(-302,11),
TO_SIGNED(-345,11),
TO_SIGNED(-386,11),
TO_SIGNED(-425,11),
TO_SIGNED(-463,11),
TO_SIGNED(-499,11),
TO_SIGNED(-533,11),
TO_SIGNED(-565,11),
TO_SIGNED(-595,11),
TO_SIGNED(-622,11),
TO_SIGNED(-647,11),
TO_SIGNED(-670,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-721,11),
TO_SIGNED(-733,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-720,11),
TO_SIGNED(-705,11),
TO_SIGNED(-688,11),
TO_SIGNED(-667,11),
TO_SIGNED(-645,11),
TO_SIGNED(-619,11),
TO_SIGNED(-592,11),
TO_SIGNED(-562,11),
TO_SIGNED(-529,11),
TO_SIGNED(-495,11),
TO_SIGNED(-459,11),
TO_SIGNED(-421,11),
TO_SIGNED(-381,11),
TO_SIGNED(-340,11),
TO_SIGNED(-297,11),
TO_SIGNED(-254,11),
TO_SIGNED(-209,11),
TO_SIGNED(-163,11),
TO_SIGNED(-117,11),
TO_SIGNED(-70,11),
TO_SIGNED(-24,11),
TO_SIGNED(24,11),
TO_SIGNED(70,11),
TO_SIGNED(117,11),
TO_SIGNED(163,11),
TO_SIGNED(209,11),
TO_SIGNED(254,11),
TO_SIGNED(297,11),
TO_SIGNED(340,11),
TO_SIGNED(381,11),
TO_SIGNED(421,11),
TO_SIGNED(459,11),
TO_SIGNED(495,11),
TO_SIGNED(529,11),
TO_SIGNED(562,11),
TO_SIGNED(592,11),
TO_SIGNED(619,11),
TO_SIGNED(645,11),
TO_SIGNED(667,11),
TO_SIGNED(688,11),
TO_SIGNED(705,11),
TO_SIGNED(720,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(733,11),
TO_SIGNED(721,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(670,11),
TO_SIGNED(647,11),
TO_SIGNED(622,11),
TO_SIGNED(595,11),
TO_SIGNED(565,11),
TO_SIGNED(533,11),
TO_SIGNED(499,11),
TO_SIGNED(463,11),
TO_SIGNED(425,11),
TO_SIGNED(386,11),
TO_SIGNED(345,11),
TO_SIGNED(302,11),
TO_SIGNED(259,11),
TO_SIGNED(214,11),
TO_SIGNED(168,11),
TO_SIGNED(122,11),
TO_SIGNED(76,11),
TO_SIGNED(29,11),
TO_SIGNED(-18,11),
TO_SIGNED(-65,11),
TO_SIGNED(-112,11),
TO_SIGNED(-158,11),
TO_SIGNED(-204,11),
TO_SIGNED(-248,11),
TO_SIGNED(-292,11),
TO_SIGNED(-335,11),
TO_SIGNED(-376,11),
TO_SIGNED(-416,11),
TO_SIGNED(-455,11),
TO_SIGNED(-491,11),
TO_SIGNED(-526,11),
TO_SIGNED(-558,11),
TO_SIGNED(-588,11),
TO_SIGNED(-616,11),
TO_SIGNED(-642,11),
TO_SIGNED(-665,11),
TO_SIGNED(-685,11),
TO_SIGNED(-703,11),
TO_SIGNED(-718,11),
TO_SIGNED(-730,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-692,11),
TO_SIGNED(-672,11),
TO_SIGNED(-650,11),
TO_SIGNED(-625,11),
TO_SIGNED(-598,11),
TO_SIGNED(-569,11),
TO_SIGNED(-537,11),
TO_SIGNED(-503,11),
TO_SIGNED(-467,11),
TO_SIGNED(-430,11),
TO_SIGNED(-390,11),
TO_SIGNED(-349,11),
TO_SIGNED(-307,11),
TO_SIGNED(-264,11),
TO_SIGNED(-219,11),
TO_SIGNED(-174,11),
TO_SIGNED(-128,11),
TO_SIGNED(-81,11),
TO_SIGNED(-34,11),
TO_SIGNED(13,11),
TO_SIGNED(60,11),
TO_SIGNED(106,11),
TO_SIGNED(153,11),
TO_SIGNED(198,11),
TO_SIGNED(243,11),
TO_SIGNED(287,11),
TO_SIGNED(330,11),
TO_SIGNED(372,11),
TO_SIGNED(412,11),
TO_SIGNED(450,11),
TO_SIGNED(487,11),
TO_SIGNED(522,11),
TO_SIGNED(554,11),
TO_SIGNED(585,11),
TO_SIGNED(613,11),
TO_SIGNED(639,11),
TO_SIGNED(662,11),
TO_SIGNED(683,11),
TO_SIGNED(701,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(724,11),
TO_SIGNED(710,11),
TO_SIGNED(694,11),
TO_SIGNED(675,11),
TO_SIGNED(653,11),
TO_SIGNED(628,11),
TO_SIGNED(601,11),
TO_SIGNED(572,11),
TO_SIGNED(541,11),
TO_SIGNED(507,11),
TO_SIGNED(471,11),
TO_SIGNED(434,11),
TO_SIGNED(395,11),
TO_SIGNED(354,11),
TO_SIGNED(312,11),
TO_SIGNED(269,11),
TO_SIGNED(224,11),
TO_SIGNED(179,11),
TO_SIGNED(133,11),
TO_SIGNED(86,11),
TO_SIGNED(40,11),
TO_SIGNED(-7,11),
TO_SIGNED(-54,11),
TO_SIGNED(-101,11),
TO_SIGNED(-148,11),
TO_SIGNED(-193,11),
TO_SIGNED(-238,11),
TO_SIGNED(-282,11),
TO_SIGNED(-325,11),
TO_SIGNED(-367,11),
TO_SIGNED(-407,11),
TO_SIGNED(-446,11),
TO_SIGNED(-483,11),
TO_SIGNED(-518,11),
TO_SIGNED(-551,11),
TO_SIGNED(-582,11),
TO_SIGNED(-610,11),
TO_SIGNED(-636,11),
TO_SIGNED(-660,11),
TO_SIGNED(-681,11),
TO_SIGNED(-699,11),
TO_SIGNED(-715,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-736,11),
TO_SIGNED(-725,11),
TO_SIGNED(-712,11),
TO_SIGNED(-696,11),
TO_SIGNED(-677,11),
TO_SIGNED(-655,11),
TO_SIGNED(-631,11),
TO_SIGNED(-605,11),
TO_SIGNED(-576,11),
TO_SIGNED(-544,11),
TO_SIGNED(-511,11),
TO_SIGNED(-476,11),
TO_SIGNED(-438,11),
TO_SIGNED(-399,11),
TO_SIGNED(-359,11),
TO_SIGNED(-317,11),
TO_SIGNED(-274,11),
TO_SIGNED(-229,11),
TO_SIGNED(-184,11),
TO_SIGNED(-138,11),
TO_SIGNED(-92,11),
TO_SIGNED(-45,11),
TO_SIGNED(2,11),
TO_SIGNED(49,11),
TO_SIGNED(96,11),
TO_SIGNED(142,11),
TO_SIGNED(188,11),
TO_SIGNED(233,11),
TO_SIGNED(277,11),
TO_SIGNED(321,11),
TO_SIGNED(362,11),
TO_SIGNED(403,11),
TO_SIGNED(442,11),
TO_SIGNED(479,11),
TO_SIGNED(514,11),
TO_SIGNED(547,11),
TO_SIGNED(578,11),
TO_SIGNED(607,11),
TO_SIGNED(633,11),
TO_SIGNED(657,11),
TO_SIGNED(679,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(698,11),
TO_SIGNED(679,11),
TO_SIGNED(658,11),
TO_SIGNED(634,11),
TO_SIGNED(608,11),
TO_SIGNED(579,11),
TO_SIGNED(548,11),
TO_SIGNED(515,11),
TO_SIGNED(480,11),
TO_SIGNED(443,11),
TO_SIGNED(404,11),
TO_SIGNED(363,11),
TO_SIGNED(322,11),
TO_SIGNED(278,11),
TO_SIGNED(234,11),
TO_SIGNED(189,11),
TO_SIGNED(143,11),
TO_SIGNED(97,11),
TO_SIGNED(50,11),
TO_SIGNED(3,11),
TO_SIGNED(-44,11),
TO_SIGNED(-91,11),
TO_SIGNED(-137,11),
TO_SIGNED(-183,11),
TO_SIGNED(-228,11),
TO_SIGNED(-273,11),
TO_SIGNED(-316,11),
TO_SIGNED(-358,11),
TO_SIGNED(-398,11),
TO_SIGNED(-437,11),
TO_SIGNED(-475,11),
TO_SIGNED(-510,11),
TO_SIGNED(-544,11),
TO_SIGNED(-575,11),
TO_SIGNED(-604,11),
TO_SIGNED(-631,11),
TO_SIGNED(-655,11),
TO_SIGNED(-676,11),
TO_SIGNED(-695,11),
TO_SIGNED(-712,11),
TO_SIGNED(-725,11),
TO_SIGNED(-736,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-715,11),
TO_SIGNED(-700,11),
TO_SIGNED(-681,11),
TO_SIGNED(-660,11),
TO_SIGNED(-637,11),
TO_SIGNED(-611,11),
TO_SIGNED(-582,11),
TO_SIGNED(-552,11),
TO_SIGNED(-519,11),
TO_SIGNED(-484,11),
TO_SIGNED(-447,11),
TO_SIGNED(-408,11),
TO_SIGNED(-368,11),
TO_SIGNED(-326,11),
TO_SIGNED(-283,11),
TO_SIGNED(-239,11),
TO_SIGNED(-194,11),
TO_SIGNED(-149,11),
TO_SIGNED(-102,11),
TO_SIGNED(-56,11),
TO_SIGNED(-9,11),
TO_SIGNED(38,11),
TO_SIGNED(85,11),
TO_SIGNED(132,11),
TO_SIGNED(178,11),
TO_SIGNED(223,11),
TO_SIGNED(268,11),
TO_SIGNED(311,11),
TO_SIGNED(353,11),
TO_SIGNED(394,11),
TO_SIGNED(433,11),
TO_SIGNED(471,11),
TO_SIGNED(506,11),
TO_SIGNED(540,11),
TO_SIGNED(571,11),
TO_SIGNED(601,11),
TO_SIGNED(628,11),
TO_SIGNED(652,11),
TO_SIGNED(674,11),
TO_SIGNED(693,11),
TO_SIGNED(710,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(739,11),
TO_SIGNED(729,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(684,11),
TO_SIGNED(663,11),
TO_SIGNED(640,11),
TO_SIGNED(614,11),
TO_SIGNED(586,11),
TO_SIGNED(555,11),
TO_SIGNED(523,11),
TO_SIGNED(488,11),
TO_SIGNED(451,11),
TO_SIGNED(413,11),
TO_SIGNED(373,11),
TO_SIGNED(331,11),
TO_SIGNED(288,11),
TO_SIGNED(244,11),
TO_SIGNED(200,11),
TO_SIGNED(154,11),
TO_SIGNED(108,11),
TO_SIGNED(61,11),
TO_SIGNED(14,11),
TO_SIGNED(-33,11),
TO_SIGNED(-80,11),
TO_SIGNED(-127,11),
TO_SIGNED(-173,11),
TO_SIGNED(-218,11),
TO_SIGNED(-263,11),
TO_SIGNED(-306,11),
TO_SIGNED(-348,11),
TO_SIGNED(-389,11),
TO_SIGNED(-429,11),
TO_SIGNED(-466,11),
TO_SIGNED(-502,11),
TO_SIGNED(-536,11),
TO_SIGNED(-568,11),
TO_SIGNED(-598,11),
TO_SIGNED(-625,11),
TO_SIGNED(-650,11),
TO_SIGNED(-672,11),
TO_SIGNED(-691,11),
TO_SIGNED(-708,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-686,11),
TO_SIGNED(-665,11),
TO_SIGNED(-642,11),
TO_SIGNED(-617,11),
TO_SIGNED(-589,11),
TO_SIGNED(-559,11),
TO_SIGNED(-526,11),
TO_SIGNED(-492,11),
TO_SIGNED(-455,11),
TO_SIGNED(-417,11),
TO_SIGNED(-377,11),
TO_SIGNED(-336,11),
TO_SIGNED(-293,11),
TO_SIGNED(-249,11),
TO_SIGNED(-205,11),
TO_SIGNED(-159,11),
TO_SIGNED(-113,11),
TO_SIGNED(-66,11),
TO_SIGNED(-19,11),
TO_SIGNED(28,11),
TO_SIGNED(75,11),
TO_SIGNED(121,11),
TO_SIGNED(167,11),
TO_SIGNED(213,11),
TO_SIGNED(258,11),
TO_SIGNED(301,11),
TO_SIGNED(344,11),
TO_SIGNED(385,11),
TO_SIGNED(424,11),
TO_SIGNED(462,11),
TO_SIGNED(498,11),
TO_SIGNED(532,11),
TO_SIGNED(564,11),
TO_SIGNED(594,11),
TO_SIGNED(622,11),
TO_SIGNED(647,11),
TO_SIGNED(669,11),
TO_SIGNED(689,11),
TO_SIGNED(706,11),
TO_SIGNED(721,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(720,11),
TO_SIGNED(705,11),
TO_SIGNED(688,11),
TO_SIGNED(668,11),
TO_SIGNED(645,11),
TO_SIGNED(620,11),
TO_SIGNED(592,11),
TO_SIGNED(562,11),
TO_SIGNED(530,11),
TO_SIGNED(496,11),
TO_SIGNED(460,11),
TO_SIGNED(422,11),
TO_SIGNED(382,11),
TO_SIGNED(341,11),
TO_SIGNED(298,11),
TO_SIGNED(255,11),
TO_SIGNED(210,11),
TO_SIGNED(164,11),
TO_SIGNED(118,11),
TO_SIGNED(71,11),
TO_SIGNED(25,11),
TO_SIGNED(-22,11),
TO_SIGNED(-69,11),
TO_SIGNED(-116,11),
TO_SIGNED(-162,11),
TO_SIGNED(-208,11),
TO_SIGNED(-252,11),
TO_SIGNED(-296,11),
TO_SIGNED(-339,11),
TO_SIGNED(-380,11),
TO_SIGNED(-420,11),
TO_SIGNED(-458,11),
TO_SIGNED(-494,11),
TO_SIGNED(-529,11),
TO_SIGNED(-561,11),
TO_SIGNED(-591,11),
TO_SIGNED(-619,11),
TO_SIGNED(-644,11),
TO_SIGNED(-667,11),
TO_SIGNED(-687,11),
TO_SIGNED(-705,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-733,11),
TO_SIGNED(-721,11),
TO_SIGNED(-707,11),
TO_SIGNED(-690,11),
TO_SIGNED(-670,11),
TO_SIGNED(-648,11),
TO_SIGNED(-623,11),
TO_SIGNED(-596,11),
TO_SIGNED(-566,11),
TO_SIGNED(-534,11),
TO_SIGNED(-500,11),
TO_SIGNED(-464,11),
TO_SIGNED(-426,11),
TO_SIGNED(-387,11),
TO_SIGNED(-345,11),
TO_SIGNED(-303,11),
TO_SIGNED(-260,11),
TO_SIGNED(-215,11),
TO_SIGNED(-169,11),
TO_SIGNED(-123,11),
TO_SIGNED(-77,11),
TO_SIGNED(-30,11),
TO_SIGNED(17,11),
TO_SIGNED(64,11),
TO_SIGNED(111,11),
TO_SIGNED(157,11),
TO_SIGNED(203,11),
TO_SIGNED(247,11),
TO_SIGNED(291,11),
TO_SIGNED(334,11),
TO_SIGNED(375,11),
TO_SIGNED(415,11),
TO_SIGNED(454,11),
TO_SIGNED(490,11),
TO_SIGNED(525,11),
TO_SIGNED(557,11),
TO_SIGNED(588,11),
TO_SIGNED(616,11),
TO_SIGNED(641,11),
TO_SIGNED(664,11),
TO_SIGNED(685,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(709,11),
TO_SIGNED(692,11),
TO_SIGNED(673,11),
TO_SIGNED(651,11),
TO_SIGNED(626,11),
TO_SIGNED(599,11),
TO_SIGNED(569,11),
TO_SIGNED(538,11),
TO_SIGNED(504,11),
TO_SIGNED(468,11),
TO_SIGNED(430,11),
TO_SIGNED(391,11),
TO_SIGNED(350,11),
TO_SIGNED(308,11),
TO_SIGNED(265,11),
TO_SIGNED(220,11),
TO_SIGNED(175,11),
TO_SIGNED(129,11),
TO_SIGNED(82,11),
TO_SIGNED(35,11),
TO_SIGNED(-12,11),
TO_SIGNED(-59,11),
TO_SIGNED(-105,11),
TO_SIGNED(-152,11),
TO_SIGNED(-197,11),
TO_SIGNED(-242,11),
TO_SIGNED(-286,11),
TO_SIGNED(-329,11),
TO_SIGNED(-371,11),
TO_SIGNED(-411,11),
TO_SIGNED(-449,11),
TO_SIGNED(-486,11),
TO_SIGNED(-521,11),
TO_SIGNED(-554,11),
TO_SIGNED(-584,11),
TO_SIGNED(-613,11),
TO_SIGNED(-639,11),
TO_SIGNED(-662,11),
TO_SIGNED(-683,11),
TO_SIGNED(-701,11),
TO_SIGNED(-716,11),
TO_SIGNED(-729,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-711,11),
TO_SIGNED(-694,11),
TO_SIGNED(-675,11),
TO_SIGNED(-653,11),
TO_SIGNED(-629,11),
TO_SIGNED(-602,11),
TO_SIGNED(-573,11),
TO_SIGNED(-541,11),
TO_SIGNED(-508,11),
TO_SIGNED(-472,11),
TO_SIGNED(-435,11),
TO_SIGNED(-396,11),
TO_SIGNED(-355,11),
TO_SIGNED(-313,11),
TO_SIGNED(-270,11),
TO_SIGNED(-225,11),
TO_SIGNED(-180,11),
TO_SIGNED(-134,11),
TO_SIGNED(-87,11),
TO_SIGNED(-41,11),
TO_SIGNED(6,11),
TO_SIGNED(53,11),
TO_SIGNED(100,11),
TO_SIGNED(147,11),
TO_SIGNED(192,11),
TO_SIGNED(237,11),
TO_SIGNED(281,11),
TO_SIGNED(324,11),
TO_SIGNED(366,11),
TO_SIGNED(406,11),
TO_SIGNED(445,11),
TO_SIGNED(482,11),
TO_SIGNED(517,11),
TO_SIGNED(550,11),
TO_SIGNED(581,11),
TO_SIGNED(610,11),
TO_SIGNED(636,11),
TO_SIGNED(659,11),
TO_SIGNED(681,11),
TO_SIGNED(699,11),
TO_SIGNED(715,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(712,11),
TO_SIGNED(696,11),
TO_SIGNED(677,11),
TO_SIGNED(656,11),
TO_SIGNED(632,11),
TO_SIGNED(605,11),
TO_SIGNED(576,11),
TO_SIGNED(545,11),
TO_SIGNED(512,11),
TO_SIGNED(476,11),
TO_SIGNED(439,11),
TO_SIGNED(400,11),
TO_SIGNED(360,11),
TO_SIGNED(318,11),
TO_SIGNED(275,11),
TO_SIGNED(230,11),
TO_SIGNED(185,11),
TO_SIGNED(139,11),
TO_SIGNED(93,11),
TO_SIGNED(46,11),
TO_SIGNED(-1,11),
TO_SIGNED(-48,11),
TO_SIGNED(-95,11),
TO_SIGNED(-141,11),
TO_SIGNED(-187,11),
TO_SIGNED(-232,11),
TO_SIGNED(-276,11),
TO_SIGNED(-320,11),
TO_SIGNED(-362,11),
TO_SIGNED(-402,11),
TO_SIGNED(-441,11),
TO_SIGNED(-478,11),
TO_SIGNED(-513,11),
TO_SIGNED(-547,11),
TO_SIGNED(-578,11),
TO_SIGNED(-606,11),
TO_SIGNED(-633,11),
TO_SIGNED(-657,11),
TO_SIGNED(-678,11),
TO_SIGNED(-697,11),
TO_SIGNED(-713,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-714,11),
TO_SIGNED(-698,11),
TO_SIGNED(-680,11),
TO_SIGNED(-658,11),
TO_SIGNED(-635,11),
TO_SIGNED(-608,11),
TO_SIGNED(-580,11),
TO_SIGNED(-549,11),
TO_SIGNED(-516,11),
TO_SIGNED(-480,11),
TO_SIGNED(-443,11),
TO_SIGNED(-405,11),
TO_SIGNED(-364,11),
TO_SIGNED(-323,11),
TO_SIGNED(-279,11),
TO_SIGNED(-235,11),
TO_SIGNED(-190,11),
TO_SIGNED(-144,11),
TO_SIGNED(-98,11),
TO_SIGNED(-51,11),
TO_SIGNED(-4,11),
TO_SIGNED(43,11),
TO_SIGNED(90,11),
TO_SIGNED(136,11),
TO_SIGNED(182,11),
TO_SIGNED(227,11),
TO_SIGNED(272,11),
TO_SIGNED(315,11),
TO_SIGNED(357,11),
TO_SIGNED(397,11),
TO_SIGNED(437,11),
TO_SIGNED(474,11),
TO_SIGNED(509,11),
TO_SIGNED(543,11),
TO_SIGNED(574,11),
TO_SIGNED(603,11),
TO_SIGNED(630,11),
TO_SIGNED(654,11),
TO_SIGNED(676,11),
TO_SIGNED(695,11),
TO_SIGNED(711,11),
TO_SIGNED(725,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(716,11),
TO_SIGNED(700,11),
TO_SIGNED(682,11),
TO_SIGNED(661,11),
TO_SIGNED(637,11),
TO_SIGNED(611,11),
TO_SIGNED(583,11),
TO_SIGNED(552,11),
TO_SIGNED(519,11),
TO_SIGNED(485,11),
TO_SIGNED(448,11),
TO_SIGNED(409,11),
TO_SIGNED(369,11),
TO_SIGNED(327,11),
TO_SIGNED(284,11),
TO_SIGNED(240,11),
TO_SIGNED(195,11),
TO_SIGNED(150,11),
TO_SIGNED(103,11),
TO_SIGNED(57,11),
TO_SIGNED(10,11),
TO_SIGNED(-37,11),
TO_SIGNED(-84,11),
TO_SIGNED(-131,11),
TO_SIGNED(-177,11),
TO_SIGNED(-222,11),
TO_SIGNED(-267,11),
TO_SIGNED(-310,11),
TO_SIGNED(-352,11),
TO_SIGNED(-393,11),
TO_SIGNED(-432,11),
TO_SIGNED(-470,11),
TO_SIGNED(-505,11),
TO_SIGNED(-539,11),
TO_SIGNED(-571,11),
TO_SIGNED(-600,11),
TO_SIGNED(-627,11),
TO_SIGNED(-652,11),
TO_SIGNED(-674,11),
TO_SIGNED(-693,11),
TO_SIGNED(-710,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-702,11),
TO_SIGNED(-684,11),
TO_SIGNED(-663,11),
TO_SIGNED(-640,11),
TO_SIGNED(-615,11),
TO_SIGNED(-586,11),
TO_SIGNED(-556,11),
TO_SIGNED(-523,11),
TO_SIGNED(-489,11),
TO_SIGNED(-452,11),
TO_SIGNED(-414,11),
TO_SIGNED(-374,11),
TO_SIGNED(-332,11),
TO_SIGNED(-289,11),
TO_SIGNED(-245,11),
TO_SIGNED(-201,11),
TO_SIGNED(-155,11),
TO_SIGNED(-109,11),
TO_SIGNED(-62,11),
TO_SIGNED(-15,11),
TO_SIGNED(32,11),
TO_SIGNED(79,11),
TO_SIGNED(125,11),
TO_SIGNED(172,11),
TO_SIGNED(217,11),
TO_SIGNED(262,11),
TO_SIGNED(305,11),
TO_SIGNED(347,11),
TO_SIGNED(388,11),
TO_SIGNED(428,11),
TO_SIGNED(466,11),
TO_SIGNED(501,11),
TO_SIGNED(535,11),
TO_SIGNED(567,11),
TO_SIGNED(597,11),
TO_SIGNED(624,11),
TO_SIGNED(649,11),
TO_SIGNED(671,11),
TO_SIGNED(691,11),
TO_SIGNED(708,11),
TO_SIGNED(722,11),
TO_SIGNED(733,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(704,11),
TO_SIGNED(686,11),
TO_SIGNED(666,11),
TO_SIGNED(643,11),
TO_SIGNED(618,11),
TO_SIGNED(590,11),
TO_SIGNED(559,11),
TO_SIGNED(527,11),
TO_SIGNED(493,11),
TO_SIGNED(456,11),
TO_SIGNED(418,11),
TO_SIGNED(378,11),
TO_SIGNED(337,11),
TO_SIGNED(294,11),
TO_SIGNED(250,11),
TO_SIGNED(206,11),
TO_SIGNED(160,11),
TO_SIGNED(114,11),
TO_SIGNED(67,11),
TO_SIGNED(20,11),
TO_SIGNED(-27,11),
TO_SIGNED(-74,11),
TO_SIGNED(-120,11),
TO_SIGNED(-166,11),
TO_SIGNED(-212,11),
TO_SIGNED(-257,11),
TO_SIGNED(-300,11),
TO_SIGNED(-343,11),
TO_SIGNED(-384,11),
TO_SIGNED(-423,11),
TO_SIGNED(-461,11),
TO_SIGNED(-497,11),
TO_SIGNED(-532,11),
TO_SIGNED(-564,11),
TO_SIGNED(-594,11),
TO_SIGNED(-621,11),
TO_SIGNED(-646,11),
TO_SIGNED(-669,11),
TO_SIGNED(-689,11),
TO_SIGNED(-706,11),
TO_SIGNED(-721,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-720,11),
TO_SIGNED(-706,11),
TO_SIGNED(-688,11),
TO_SIGNED(-668,11),
TO_SIGNED(-646,11),
TO_SIGNED(-621,11),
TO_SIGNED(-593,11),
TO_SIGNED(-563,11),
TO_SIGNED(-531,11),
TO_SIGNED(-497,11),
TO_SIGNED(-460,11),
TO_SIGNED(-422,11),
TO_SIGNED(-383,11),
TO_SIGNED(-342,11),
TO_SIGNED(-299,11),
TO_SIGNED(-256,11),
TO_SIGNED(-211,11),
TO_SIGNED(-165,11),
TO_SIGNED(-119,11),
TO_SIGNED(-73,11),
TO_SIGNED(-26,11),
TO_SIGNED(21,11),
TO_SIGNED(68,11),
TO_SIGNED(115,11),
TO_SIGNED(161,11),
TO_SIGNED(207,11),
TO_SIGNED(251,11),
TO_SIGNED(295,11),
TO_SIGNED(338,11),
TO_SIGNED(379,11),
TO_SIGNED(419,11),
TO_SIGNED(457,11),
TO_SIGNED(493,11),
TO_SIGNED(528,11),
TO_SIGNED(560,11),
TO_SIGNED(590,11),
TO_SIGNED(618,11),
TO_SIGNED(644,11),
TO_SIGNED(666,11),
TO_SIGNED(687,11),
TO_SIGNED(704,11),
TO_SIGNED(719,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(671,11),
TO_SIGNED(648,11),
TO_SIGNED(624,11),
TO_SIGNED(596,11),
TO_SIGNED(567,11),
TO_SIGNED(535,11),
TO_SIGNED(501,11),
TO_SIGNED(465,11),
TO_SIGNED(427,11),
TO_SIGNED(387,11),
TO_SIGNED(346,11),
TO_SIGNED(304,11),
TO_SIGNED(261,11),
TO_SIGNED(216,11),
TO_SIGNED(171,11),
TO_SIGNED(124,11),
TO_SIGNED(78,11),
TO_SIGNED(31,11),
TO_SIGNED(-16,11),
TO_SIGNED(-63,11),
TO_SIGNED(-110,11),
TO_SIGNED(-156,11),
TO_SIGNED(-202,11),
TO_SIGNED(-246,11),
TO_SIGNED(-290,11),
TO_SIGNED(-333,11),
TO_SIGNED(-375,11),
TO_SIGNED(-415,11),
TO_SIGNED(-453,11),
TO_SIGNED(-489,11),
TO_SIGNED(-524,11),
TO_SIGNED(-557,11),
TO_SIGNED(-587,11),
TO_SIGNED(-615,11),
TO_SIGNED(-641,11),
TO_SIGNED(-664,11),
TO_SIGNED(-685,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-730,11),
TO_SIGNED(-739,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-693,11),
TO_SIGNED(-673,11),
TO_SIGNED(-651,11),
TO_SIGNED(-627,11),
TO_SIGNED(-599,11),
TO_SIGNED(-570,11),
TO_SIGNED(-538,11),
TO_SIGNED(-505,11),
TO_SIGNED(-469,11),
TO_SIGNED(-431,11),
TO_SIGNED(-392,11),
TO_SIGNED(-351,11),
TO_SIGNED(-309,11),
TO_SIGNED(-266,11),
TO_SIGNED(-221,11),
TO_SIGNED(-176,11),
TO_SIGNED(-130,11),
TO_SIGNED(-83,11),
TO_SIGNED(-36,11),
TO_SIGNED(11,11),
TO_SIGNED(58,11),
TO_SIGNED(104,11),
TO_SIGNED(151,11),
TO_SIGNED(196,11),
TO_SIGNED(241,11),
TO_SIGNED(285,11),
TO_SIGNED(328,11),
TO_SIGNED(370,11),
TO_SIGNED(410,11),
TO_SIGNED(449,11),
TO_SIGNED(485,11),
TO_SIGNED(520,11),
TO_SIGNED(553,11),
TO_SIGNED(584,11),
TO_SIGNED(612,11),
TO_SIGNED(638,11),
TO_SIGNED(661,11),
TO_SIGNED(682,11),
TO_SIGNED(700,11),
TO_SIGNED(716,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(725,11),
TO_SIGNED(711,11),
TO_SIGNED(695,11),
TO_SIGNED(675,11),
TO_SIGNED(654,11),
TO_SIGNED(629,11),
TO_SIGNED(603,11),
TO_SIGNED(574,11),
TO_SIGNED(542,11),
TO_SIGNED(509,11),
TO_SIGNED(473,11),
TO_SIGNED(436,11),
TO_SIGNED(397,11),
TO_SIGNED(356,11),
TO_SIGNED(314,11),
TO_SIGNED(271,11),
TO_SIGNED(226,11),
TO_SIGNED(181,11),
TO_SIGNED(135,11),
TO_SIGNED(88,11),
TO_SIGNED(42,11),
TO_SIGNED(-5,11),
TO_SIGNED(-52,11),
TO_SIGNED(-99,11),
TO_SIGNED(-145,11),
TO_SIGNED(-191,11),
TO_SIGNED(-236,11),
TO_SIGNED(-280,11),
TO_SIGNED(-323,11),
TO_SIGNED(-365,11),
TO_SIGNED(-406,11),
TO_SIGNED(-444,11),
TO_SIGNED(-481,11),
TO_SIGNED(-516,11),
TO_SIGNED(-549,11),
TO_SIGNED(-580,11),
TO_SIGNED(-609,11),
TO_SIGNED(-635,11),
TO_SIGNED(-659,11),
TO_SIGNED(-680,11),
TO_SIGNED(-699,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-736,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-678,11),
TO_SIGNED(-656,11),
TO_SIGNED(-632,11),
TO_SIGNED(-606,11),
TO_SIGNED(-577,11),
TO_SIGNED(-546,11),
TO_SIGNED(-512,11),
TO_SIGNED(-477,11),
TO_SIGNED(-440,11),
TO_SIGNED(-401,11),
TO_SIGNED(-361,11),
TO_SIGNED(-319,11),
TO_SIGNED(-275,11),
TO_SIGNED(-231,11),
TO_SIGNED(-186,11),
TO_SIGNED(-140,11),
TO_SIGNED(-94,11),
TO_SIGNED(-47,11),
TO_SIGNED(0,11),
TO_SIGNED(47,11),
TO_SIGNED(94,11),
TO_SIGNED(140,11),
TO_SIGNED(186,11),
TO_SIGNED(231,11),
TO_SIGNED(275,11),
TO_SIGNED(319,11),
TO_SIGNED(361,11),
TO_SIGNED(401,11),
TO_SIGNED(440,11),
TO_SIGNED(477,11),
TO_SIGNED(512,11),
TO_SIGNED(546,11),
TO_SIGNED(577,11),
TO_SIGNED(606,11),
TO_SIGNED(632,11),
TO_SIGNED(656,11),
TO_SIGNED(678,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(736,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(699,11),
TO_SIGNED(680,11),
TO_SIGNED(659,11),
TO_SIGNED(635,11),
TO_SIGNED(609,11),
TO_SIGNED(580,11),
TO_SIGNED(549,11),
TO_SIGNED(516,11),
TO_SIGNED(481,11),
TO_SIGNED(444,11),
TO_SIGNED(406,11),
TO_SIGNED(365,11),
TO_SIGNED(323,11),
TO_SIGNED(280,11),
TO_SIGNED(236,11),
TO_SIGNED(191,11),
TO_SIGNED(145,11),
TO_SIGNED(99,11),
TO_SIGNED(52,11),
TO_SIGNED(5,11),
TO_SIGNED(-42,11),
TO_SIGNED(-88,11),
TO_SIGNED(-135,11),
TO_SIGNED(-181,11),
TO_SIGNED(-226,11),
TO_SIGNED(-271,11),
TO_SIGNED(-314,11),
TO_SIGNED(-356,11),
TO_SIGNED(-397,11),
TO_SIGNED(-436,11),
TO_SIGNED(-473,11),
TO_SIGNED(-509,11),
TO_SIGNED(-542,11),
TO_SIGNED(-574,11),
TO_SIGNED(-603,11),
TO_SIGNED(-629,11),
TO_SIGNED(-654,11),
TO_SIGNED(-675,11),
TO_SIGNED(-695,11),
TO_SIGNED(-711,11),
TO_SIGNED(-725,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-716,11),
TO_SIGNED(-700,11),
TO_SIGNED(-682,11),
TO_SIGNED(-661,11),
TO_SIGNED(-638,11),
TO_SIGNED(-612,11),
TO_SIGNED(-584,11),
TO_SIGNED(-553,11),
TO_SIGNED(-520,11),
TO_SIGNED(-485,11),
TO_SIGNED(-449,11),
TO_SIGNED(-410,11),
TO_SIGNED(-370,11),
TO_SIGNED(-328,11),
TO_SIGNED(-285,11),
TO_SIGNED(-241,11),
TO_SIGNED(-196,11),
TO_SIGNED(-151,11),
TO_SIGNED(-104,11),
TO_SIGNED(-58,11),
TO_SIGNED(-11,11),
TO_SIGNED(36,11),
TO_SIGNED(83,11),
TO_SIGNED(130,11),
TO_SIGNED(176,11),
TO_SIGNED(221,11),
TO_SIGNED(266,11),
TO_SIGNED(309,11),
TO_SIGNED(351,11),
TO_SIGNED(392,11),
TO_SIGNED(431,11),
TO_SIGNED(469,11),
TO_SIGNED(505,11),
TO_SIGNED(538,11),
TO_SIGNED(570,11),
TO_SIGNED(599,11),
TO_SIGNED(627,11),
TO_SIGNED(651,11),
TO_SIGNED(673,11),
TO_SIGNED(693,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(739,11),
TO_SIGNED(730,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(685,11),
TO_SIGNED(664,11),
TO_SIGNED(641,11),
TO_SIGNED(615,11),
TO_SIGNED(587,11),
TO_SIGNED(557,11),
TO_SIGNED(524,11),
TO_SIGNED(489,11),
TO_SIGNED(453,11),
TO_SIGNED(415,11),
TO_SIGNED(375,11),
TO_SIGNED(333,11),
TO_SIGNED(290,11),
TO_SIGNED(246,11),
TO_SIGNED(202,11),
TO_SIGNED(156,11),
TO_SIGNED(110,11),
TO_SIGNED(63,11),
TO_SIGNED(16,11),
TO_SIGNED(-31,11),
TO_SIGNED(-78,11),
TO_SIGNED(-124,11),
TO_SIGNED(-171,11),
TO_SIGNED(-216,11),
TO_SIGNED(-261,11),
TO_SIGNED(-304,11),
TO_SIGNED(-346,11),
TO_SIGNED(-387,11),
TO_SIGNED(-427,11),
TO_SIGNED(-465,11),
TO_SIGNED(-501,11),
TO_SIGNED(-535,11),
TO_SIGNED(-567,11),
TO_SIGNED(-596,11),
TO_SIGNED(-624,11),
TO_SIGNED(-648,11),
TO_SIGNED(-671,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-719,11),
TO_SIGNED(-704,11),
TO_SIGNED(-687,11),
TO_SIGNED(-666,11),
TO_SIGNED(-644,11),
TO_SIGNED(-618,11),
TO_SIGNED(-590,11),
TO_SIGNED(-560,11),
TO_SIGNED(-528,11),
TO_SIGNED(-493,11),
TO_SIGNED(-457,11),
TO_SIGNED(-419,11),
TO_SIGNED(-379,11),
TO_SIGNED(-338,11),
TO_SIGNED(-295,11),
TO_SIGNED(-251,11),
TO_SIGNED(-207,11),
TO_SIGNED(-161,11),
TO_SIGNED(-115,11),
TO_SIGNED(-68,11),
TO_SIGNED(-21,11),
TO_SIGNED(26,11),
TO_SIGNED(73,11),
TO_SIGNED(119,11),
TO_SIGNED(165,11),
TO_SIGNED(211,11),
TO_SIGNED(256,11),
TO_SIGNED(299,11),
TO_SIGNED(342,11),
TO_SIGNED(383,11),
TO_SIGNED(422,11),
TO_SIGNED(460,11),
TO_SIGNED(497,11),
TO_SIGNED(531,11),
TO_SIGNED(563,11),
TO_SIGNED(593,11),
TO_SIGNED(621,11),
TO_SIGNED(646,11),
TO_SIGNED(668,11),
TO_SIGNED(688,11),
TO_SIGNED(706,11),
TO_SIGNED(720,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(721,11),
TO_SIGNED(706,11),
TO_SIGNED(689,11),
TO_SIGNED(669,11),
TO_SIGNED(646,11),
TO_SIGNED(621,11),
TO_SIGNED(594,11),
TO_SIGNED(564,11),
TO_SIGNED(532,11),
TO_SIGNED(497,11),
TO_SIGNED(461,11),
TO_SIGNED(423,11),
TO_SIGNED(384,11),
TO_SIGNED(343,11),
TO_SIGNED(300,11),
TO_SIGNED(257,11),
TO_SIGNED(212,11),
TO_SIGNED(166,11),
TO_SIGNED(120,11),
TO_SIGNED(74,11),
TO_SIGNED(27,11),
TO_SIGNED(-20,11),
TO_SIGNED(-67,11),
TO_SIGNED(-114,11),
TO_SIGNED(-160,11),
TO_SIGNED(-206,11),
TO_SIGNED(-250,11),
TO_SIGNED(-294,11),
TO_SIGNED(-337,11),
TO_SIGNED(-378,11),
TO_SIGNED(-418,11),
TO_SIGNED(-456,11),
TO_SIGNED(-493,11),
TO_SIGNED(-527,11),
TO_SIGNED(-559,11),
TO_SIGNED(-590,11),
TO_SIGNED(-618,11),
TO_SIGNED(-643,11),
TO_SIGNED(-666,11),
TO_SIGNED(-686,11),
TO_SIGNED(-704,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-733,11),
TO_SIGNED(-722,11),
TO_SIGNED(-708,11),
TO_SIGNED(-691,11),
TO_SIGNED(-671,11),
TO_SIGNED(-649,11),
TO_SIGNED(-624,11),
TO_SIGNED(-597,11),
TO_SIGNED(-567,11),
TO_SIGNED(-535,11),
TO_SIGNED(-501,11),
TO_SIGNED(-466,11),
TO_SIGNED(-428,11),
TO_SIGNED(-388,11),
TO_SIGNED(-347,11),
TO_SIGNED(-305,11),
TO_SIGNED(-262,11),
TO_SIGNED(-217,11),
TO_SIGNED(-172,11),
TO_SIGNED(-125,11),
TO_SIGNED(-79,11),
TO_SIGNED(-32,11),
TO_SIGNED(15,11),
TO_SIGNED(62,11),
TO_SIGNED(109,11),
TO_SIGNED(155,11),
TO_SIGNED(201,11),
TO_SIGNED(245,11),
TO_SIGNED(289,11),
TO_SIGNED(332,11),
TO_SIGNED(374,11),
TO_SIGNED(414,11),
TO_SIGNED(452,11),
TO_SIGNED(489,11),
TO_SIGNED(523,11),
TO_SIGNED(556,11),
TO_SIGNED(586,11),
TO_SIGNED(615,11),
TO_SIGNED(640,11),
TO_SIGNED(663,11),
TO_SIGNED(684,11),
TO_SIGNED(702,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(710,11),
TO_SIGNED(693,11),
TO_SIGNED(674,11),
TO_SIGNED(652,11),
TO_SIGNED(627,11),
TO_SIGNED(600,11),
TO_SIGNED(571,11),
TO_SIGNED(539,11),
TO_SIGNED(505,11),
TO_SIGNED(470,11),
TO_SIGNED(432,11),
TO_SIGNED(393,11),
TO_SIGNED(352,11),
TO_SIGNED(310,11),
TO_SIGNED(267,11),
TO_SIGNED(222,11),
TO_SIGNED(177,11),
TO_SIGNED(131,11),
TO_SIGNED(84,11),
TO_SIGNED(37,11),
TO_SIGNED(-10,11),
TO_SIGNED(-57,11),
TO_SIGNED(-103,11),
TO_SIGNED(-150,11),
TO_SIGNED(-195,11),
TO_SIGNED(-240,11),
TO_SIGNED(-284,11),
TO_SIGNED(-327,11),
TO_SIGNED(-369,11),
TO_SIGNED(-409,11),
TO_SIGNED(-448,11),
TO_SIGNED(-485,11),
TO_SIGNED(-519,11),
TO_SIGNED(-552,11),
TO_SIGNED(-583,11),
TO_SIGNED(-611,11),
TO_SIGNED(-637,11),
TO_SIGNED(-661,11),
TO_SIGNED(-682,11),
TO_SIGNED(-700,11),
TO_SIGNED(-716,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-725,11),
TO_SIGNED(-711,11),
TO_SIGNED(-695,11),
TO_SIGNED(-676,11),
TO_SIGNED(-654,11),
TO_SIGNED(-630,11),
TO_SIGNED(-603,11),
TO_SIGNED(-574,11),
TO_SIGNED(-543,11),
TO_SIGNED(-509,11),
TO_SIGNED(-474,11),
TO_SIGNED(-437,11),
TO_SIGNED(-397,11),
TO_SIGNED(-357,11),
TO_SIGNED(-315,11),
TO_SIGNED(-272,11),
TO_SIGNED(-227,11),
TO_SIGNED(-182,11),
TO_SIGNED(-136,11),
TO_SIGNED(-90,11),
TO_SIGNED(-43,11),
TO_SIGNED(4,11),
TO_SIGNED(51,11),
TO_SIGNED(98,11),
TO_SIGNED(144,11),
TO_SIGNED(190,11),
TO_SIGNED(235,11),
TO_SIGNED(279,11),
TO_SIGNED(323,11),
TO_SIGNED(364,11),
TO_SIGNED(405,11),
TO_SIGNED(443,11),
TO_SIGNED(480,11),
TO_SIGNED(516,11),
TO_SIGNED(549,11),
TO_SIGNED(580,11),
TO_SIGNED(608,11),
TO_SIGNED(635,11),
TO_SIGNED(658,11),
TO_SIGNED(680,11),
TO_SIGNED(698,11),
TO_SIGNED(714,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(713,11),
TO_SIGNED(697,11),
TO_SIGNED(678,11),
TO_SIGNED(657,11),
TO_SIGNED(633,11),
TO_SIGNED(606,11),
TO_SIGNED(578,11),
TO_SIGNED(547,11),
TO_SIGNED(513,11),
TO_SIGNED(478,11),
TO_SIGNED(441,11),
TO_SIGNED(402,11),
TO_SIGNED(362,11),
TO_SIGNED(320,11),
TO_SIGNED(276,11),
TO_SIGNED(232,11),
TO_SIGNED(187,11),
TO_SIGNED(141,11),
TO_SIGNED(95,11),
TO_SIGNED(48,11),
TO_SIGNED(1,11),
TO_SIGNED(-46,11),
TO_SIGNED(-93,11),
TO_SIGNED(-139,11),
TO_SIGNED(-185,11),
TO_SIGNED(-230,11),
TO_SIGNED(-275,11),
TO_SIGNED(-318,11),
TO_SIGNED(-360,11),
TO_SIGNED(-400,11),
TO_SIGNED(-439,11),
TO_SIGNED(-476,11),
TO_SIGNED(-512,11),
TO_SIGNED(-545,11),
TO_SIGNED(-576,11),
TO_SIGNED(-605,11),
TO_SIGNED(-632,11),
TO_SIGNED(-656,11),
TO_SIGNED(-677,11),
TO_SIGNED(-696,11),
TO_SIGNED(-712,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-715,11),
TO_SIGNED(-699,11),
TO_SIGNED(-681,11),
TO_SIGNED(-659,11),
TO_SIGNED(-636,11),
TO_SIGNED(-610,11),
TO_SIGNED(-581,11),
TO_SIGNED(-550,11),
TO_SIGNED(-517,11),
TO_SIGNED(-482,11),
TO_SIGNED(-445,11),
TO_SIGNED(-406,11),
TO_SIGNED(-366,11),
TO_SIGNED(-324,11),
TO_SIGNED(-281,11),
TO_SIGNED(-237,11),
TO_SIGNED(-192,11),
TO_SIGNED(-147,11),
TO_SIGNED(-100,11),
TO_SIGNED(-53,11),
TO_SIGNED(-6,11),
TO_SIGNED(41,11),
TO_SIGNED(87,11),
TO_SIGNED(134,11),
TO_SIGNED(180,11),
TO_SIGNED(225,11),
TO_SIGNED(270,11),
TO_SIGNED(313,11),
TO_SIGNED(355,11),
TO_SIGNED(396,11),
TO_SIGNED(435,11),
TO_SIGNED(472,11),
TO_SIGNED(508,11),
TO_SIGNED(541,11),
TO_SIGNED(573,11),
TO_SIGNED(602,11),
TO_SIGNED(629,11),
TO_SIGNED(653,11),
TO_SIGNED(675,11),
TO_SIGNED(694,11),
TO_SIGNED(711,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(729,11),
TO_SIGNED(716,11),
TO_SIGNED(701,11),
TO_SIGNED(683,11),
TO_SIGNED(662,11),
TO_SIGNED(639,11),
TO_SIGNED(613,11),
TO_SIGNED(584,11),
TO_SIGNED(554,11),
TO_SIGNED(521,11),
TO_SIGNED(486,11),
TO_SIGNED(449,11),
TO_SIGNED(411,11),
TO_SIGNED(371,11),
TO_SIGNED(329,11),
TO_SIGNED(286,11),
TO_SIGNED(242,11),
TO_SIGNED(197,11),
TO_SIGNED(152,11),
TO_SIGNED(105,11),
TO_SIGNED(59,11),
TO_SIGNED(12,11),
TO_SIGNED(-35,11),
TO_SIGNED(-82,11),
TO_SIGNED(-129,11),
TO_SIGNED(-175,11),
TO_SIGNED(-220,11),
TO_SIGNED(-265,11),
TO_SIGNED(-308,11),
TO_SIGNED(-350,11),
TO_SIGNED(-391,11),
TO_SIGNED(-430,11),
TO_SIGNED(-468,11),
TO_SIGNED(-504,11),
TO_SIGNED(-538,11),
TO_SIGNED(-569,11),
TO_SIGNED(-599,11),
TO_SIGNED(-626,11),
TO_SIGNED(-651,11),
TO_SIGNED(-673,11),
TO_SIGNED(-692,11),
TO_SIGNED(-709,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-685,11),
TO_SIGNED(-664,11),
TO_SIGNED(-641,11),
TO_SIGNED(-616,11),
TO_SIGNED(-588,11),
TO_SIGNED(-557,11),
TO_SIGNED(-525,11),
TO_SIGNED(-490,11),
TO_SIGNED(-454,11),
TO_SIGNED(-415,11),
TO_SIGNED(-375,11),
TO_SIGNED(-334,11),
TO_SIGNED(-291,11),
TO_SIGNED(-247,11),
TO_SIGNED(-203,11),
TO_SIGNED(-157,11),
TO_SIGNED(-111,11),
TO_SIGNED(-64,11),
TO_SIGNED(-17,11),
TO_SIGNED(30,11),
TO_SIGNED(77,11),
TO_SIGNED(123,11),
TO_SIGNED(169,11),
TO_SIGNED(215,11),
TO_SIGNED(260,11),
TO_SIGNED(303,11),
TO_SIGNED(345,11),
TO_SIGNED(387,11),
TO_SIGNED(426,11),
TO_SIGNED(464,11),
TO_SIGNED(500,11),
TO_SIGNED(534,11),
TO_SIGNED(566,11),
TO_SIGNED(596,11),
TO_SIGNED(623,11),
TO_SIGNED(648,11),
TO_SIGNED(670,11),
TO_SIGNED(690,11),
TO_SIGNED(707,11),
TO_SIGNED(721,11),
TO_SIGNED(733,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(705,11),
TO_SIGNED(687,11),
TO_SIGNED(667,11),
TO_SIGNED(644,11),
TO_SIGNED(619,11),
TO_SIGNED(591,11),
TO_SIGNED(561,11),
TO_SIGNED(529,11),
TO_SIGNED(494,11),
TO_SIGNED(458,11),
TO_SIGNED(420,11),
TO_SIGNED(380,11),
TO_SIGNED(339,11),
TO_SIGNED(296,11),
TO_SIGNED(252,11),
TO_SIGNED(208,11),
TO_SIGNED(162,11),
TO_SIGNED(116,11),
TO_SIGNED(69,11),
TO_SIGNED(22,11),
TO_SIGNED(-25,11),
TO_SIGNED(-71,11),
TO_SIGNED(-118,11),
TO_SIGNED(-164,11),
TO_SIGNED(-210,11),
TO_SIGNED(-255,11),
TO_SIGNED(-298,11),
TO_SIGNED(-341,11),
TO_SIGNED(-382,11),
TO_SIGNED(-422,11),
TO_SIGNED(-460,11),
TO_SIGNED(-496,11),
TO_SIGNED(-530,11),
TO_SIGNED(-562,11),
TO_SIGNED(-592,11),
TO_SIGNED(-620,11),
TO_SIGNED(-645,11),
TO_SIGNED(-668,11),
TO_SIGNED(-688,11),
TO_SIGNED(-705,11),
TO_SIGNED(-720,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-721,11),
TO_SIGNED(-706,11),
TO_SIGNED(-689,11),
TO_SIGNED(-669,11),
TO_SIGNED(-647,11),
TO_SIGNED(-622,11),
TO_SIGNED(-594,11),
TO_SIGNED(-564,11),
TO_SIGNED(-532,11),
TO_SIGNED(-498,11),
TO_SIGNED(-462,11),
TO_SIGNED(-424,11),
TO_SIGNED(-385,11),
TO_SIGNED(-344,11),
TO_SIGNED(-301,11),
TO_SIGNED(-258,11),
TO_SIGNED(-213,11),
TO_SIGNED(-167,11),
TO_SIGNED(-121,11),
TO_SIGNED(-75,11),
TO_SIGNED(-28,11),
TO_SIGNED(19,11),
TO_SIGNED(66,11),
TO_SIGNED(113,11),
TO_SIGNED(159,11),
TO_SIGNED(205,11),
TO_SIGNED(249,11),
TO_SIGNED(293,11),
TO_SIGNED(336,11),
TO_SIGNED(377,11),
TO_SIGNED(417,11),
TO_SIGNED(455,11),
TO_SIGNED(492,11),
TO_SIGNED(526,11),
TO_SIGNED(559,11),
TO_SIGNED(589,11),
TO_SIGNED(617,11),
TO_SIGNED(642,11),
TO_SIGNED(665,11),
TO_SIGNED(686,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(708,11),
TO_SIGNED(691,11),
TO_SIGNED(672,11),
TO_SIGNED(650,11),
TO_SIGNED(625,11),
TO_SIGNED(598,11),
TO_SIGNED(568,11),
TO_SIGNED(536,11),
TO_SIGNED(502,11),
TO_SIGNED(466,11),
TO_SIGNED(429,11),
TO_SIGNED(389,11),
TO_SIGNED(348,11),
TO_SIGNED(306,11),
TO_SIGNED(263,11),
TO_SIGNED(218,11),
TO_SIGNED(173,11),
TO_SIGNED(127,11),
TO_SIGNED(80,11),
TO_SIGNED(33,11),
TO_SIGNED(-14,11),
TO_SIGNED(-61,11),
TO_SIGNED(-108,11),
TO_SIGNED(-154,11),
TO_SIGNED(-200,11),
TO_SIGNED(-244,11),
TO_SIGNED(-288,11),
TO_SIGNED(-331,11),
TO_SIGNED(-373,11),
TO_SIGNED(-413,11),
TO_SIGNED(-451,11),
TO_SIGNED(-488,11),
TO_SIGNED(-523,11),
TO_SIGNED(-555,11),
TO_SIGNED(-586,11),
TO_SIGNED(-614,11),
TO_SIGNED(-640,11),
TO_SIGNED(-663,11),
TO_SIGNED(-684,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-729,11),
TO_SIGNED(-739,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-710,11),
TO_SIGNED(-693,11),
TO_SIGNED(-674,11),
TO_SIGNED(-652,11),
TO_SIGNED(-628,11),
TO_SIGNED(-601,11),
TO_SIGNED(-571,11),
TO_SIGNED(-540,11),
TO_SIGNED(-506,11),
TO_SIGNED(-471,11),
TO_SIGNED(-433,11),
TO_SIGNED(-394,11),
TO_SIGNED(-353,11),
TO_SIGNED(-311,11),
TO_SIGNED(-268,11),
TO_SIGNED(-223,11),
TO_SIGNED(-178,11),
TO_SIGNED(-132,11),
TO_SIGNED(-85,11),
TO_SIGNED(-38,11),
TO_SIGNED(9,11),
TO_SIGNED(56,11),
TO_SIGNED(102,11),
TO_SIGNED(149,11),
TO_SIGNED(194,11),
TO_SIGNED(239,11),
TO_SIGNED(283,11),
TO_SIGNED(326,11),
TO_SIGNED(368,11),
TO_SIGNED(408,11),
TO_SIGNED(447,11),
TO_SIGNED(484,11),
TO_SIGNED(519,11),
TO_SIGNED(552,11),
TO_SIGNED(582,11),
TO_SIGNED(611,11),
TO_SIGNED(637,11),
TO_SIGNED(660,11),
TO_SIGNED(681,11),
TO_SIGNED(700,11),
TO_SIGNED(715,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(736,11),
TO_SIGNED(725,11),
TO_SIGNED(712,11),
TO_SIGNED(695,11),
TO_SIGNED(676,11),
TO_SIGNED(655,11),
TO_SIGNED(631,11),
TO_SIGNED(604,11),
TO_SIGNED(575,11),
TO_SIGNED(544,11),
TO_SIGNED(510,11),
TO_SIGNED(475,11),
TO_SIGNED(437,11),
TO_SIGNED(398,11),
TO_SIGNED(358,11),
TO_SIGNED(316,11),
TO_SIGNED(273,11),
TO_SIGNED(228,11),
TO_SIGNED(183,11),
TO_SIGNED(137,11),
TO_SIGNED(91,11),
TO_SIGNED(44,11),
TO_SIGNED(-3,11),
TO_SIGNED(-50,11),
TO_SIGNED(-97,11),
TO_SIGNED(-143,11),
TO_SIGNED(-189,11),
TO_SIGNED(-234,11),
TO_SIGNED(-278,11),
TO_SIGNED(-322,11),
TO_SIGNED(-363,11),
TO_SIGNED(-404,11),
TO_SIGNED(-443,11),
TO_SIGNED(-480,11),
TO_SIGNED(-515,11),
TO_SIGNED(-548,11),
TO_SIGNED(-579,11),
TO_SIGNED(-608,11),
TO_SIGNED(-634,11),
TO_SIGNED(-658,11),
TO_SIGNED(-679,11),
TO_SIGNED(-698,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-679,11),
TO_SIGNED(-657,11),
TO_SIGNED(-633,11),
TO_SIGNED(-607,11),
TO_SIGNED(-578,11),
TO_SIGNED(-547,11),
TO_SIGNED(-514,11),
TO_SIGNED(-479,11),
TO_SIGNED(-442,11),
TO_SIGNED(-403,11),
TO_SIGNED(-362,11),
TO_SIGNED(-321,11),
TO_SIGNED(-277,11),
TO_SIGNED(-233,11),
TO_SIGNED(-188,11),
TO_SIGNED(-142,11),
TO_SIGNED(-96,11),
TO_SIGNED(-49,11),
TO_SIGNED(-2,11),
TO_SIGNED(45,11),
TO_SIGNED(92,11),
TO_SIGNED(138,11),
TO_SIGNED(184,11),
TO_SIGNED(229,11),
TO_SIGNED(274,11),
TO_SIGNED(317,11),
TO_SIGNED(359,11),
TO_SIGNED(399,11),
TO_SIGNED(438,11),
TO_SIGNED(476,11),
TO_SIGNED(511,11),
TO_SIGNED(544,11),
TO_SIGNED(576,11),
TO_SIGNED(605,11),
TO_SIGNED(631,11),
TO_SIGNED(655,11),
TO_SIGNED(677,11),
TO_SIGNED(696,11),
TO_SIGNED(712,11),
TO_SIGNED(725,11),
TO_SIGNED(736,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(715,11),
TO_SIGNED(699,11),
TO_SIGNED(681,11),
TO_SIGNED(660,11),
TO_SIGNED(636,11),
TO_SIGNED(610,11),
TO_SIGNED(582,11),
TO_SIGNED(551,11),
TO_SIGNED(518,11),
TO_SIGNED(483,11),
TO_SIGNED(446,11),
TO_SIGNED(407,11),
TO_SIGNED(367,11),
TO_SIGNED(325,11),
TO_SIGNED(282,11),
TO_SIGNED(238,11),
TO_SIGNED(193,11),
TO_SIGNED(148,11),
TO_SIGNED(101,11),
TO_SIGNED(54,11),
TO_SIGNED(7,11),
TO_SIGNED(-40,11),
TO_SIGNED(-86,11),
TO_SIGNED(-133,11),
TO_SIGNED(-179,11),
TO_SIGNED(-224,11),
TO_SIGNED(-269,11),
TO_SIGNED(-312,11),
TO_SIGNED(-354,11),
TO_SIGNED(-395,11),
TO_SIGNED(-434,11),
TO_SIGNED(-471,11),
TO_SIGNED(-507,11),
TO_SIGNED(-541,11),
TO_SIGNED(-572,11),
TO_SIGNED(-601,11),
TO_SIGNED(-628,11),
TO_SIGNED(-653,11),
TO_SIGNED(-675,11),
TO_SIGNED(-694,11),
TO_SIGNED(-710,11),
TO_SIGNED(-724,11),
TO_SIGNED(-735,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-701,11),
TO_SIGNED(-683,11),
TO_SIGNED(-662,11),
TO_SIGNED(-639,11),
TO_SIGNED(-613,11),
TO_SIGNED(-585,11),
TO_SIGNED(-554,11),
TO_SIGNED(-522,11),
TO_SIGNED(-487,11),
TO_SIGNED(-450,11),
TO_SIGNED(-412,11),
TO_SIGNED(-372,11),
TO_SIGNED(-330,11),
TO_SIGNED(-287,11),
TO_SIGNED(-243,11),
TO_SIGNED(-198,11),
TO_SIGNED(-153,11),
TO_SIGNED(-106,11),
TO_SIGNED(-60,11),
TO_SIGNED(-13,11),
TO_SIGNED(34,11),
TO_SIGNED(81,11),
TO_SIGNED(128,11),
TO_SIGNED(174,11),
TO_SIGNED(219,11),
TO_SIGNED(264,11),
TO_SIGNED(307,11),
TO_SIGNED(349,11),
TO_SIGNED(390,11),
TO_SIGNED(430,11),
TO_SIGNED(467,11),
TO_SIGNED(503,11),
TO_SIGNED(537,11),
TO_SIGNED(569,11),
TO_SIGNED(598,11),
TO_SIGNED(625,11),
TO_SIGNED(650,11),
TO_SIGNED(672,11),
TO_SIGNED(692,11),
TO_SIGNED(709,11),
TO_SIGNED(723,11),
TO_SIGNED(734,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(730,11),
TO_SIGNED(718,11),
TO_SIGNED(703,11),
TO_SIGNED(685,11),
TO_SIGNED(665,11),
TO_SIGNED(642,11),
TO_SIGNED(616,11),
TO_SIGNED(588,11),
TO_SIGNED(558,11),
TO_SIGNED(526,11),
TO_SIGNED(491,11),
TO_SIGNED(455,11),
TO_SIGNED(416,11),
TO_SIGNED(376,11),
TO_SIGNED(335,11),
TO_SIGNED(292,11),
TO_SIGNED(248,11),
TO_SIGNED(204,11),
TO_SIGNED(158,11),
TO_SIGNED(112,11),
TO_SIGNED(65,11),
TO_SIGNED(18,11),
TO_SIGNED(-29,11),
TO_SIGNED(-76,11),
TO_SIGNED(-122,11),
TO_SIGNED(-168,11),
TO_SIGNED(-214,11),
TO_SIGNED(-259,11),
TO_SIGNED(-302,11),
TO_SIGNED(-345,11),
TO_SIGNED(-386,11),
TO_SIGNED(-425,11),
TO_SIGNED(-463,11),
TO_SIGNED(-499,11),
TO_SIGNED(-533,11),
TO_SIGNED(-565,11),
TO_SIGNED(-595,11),
TO_SIGNED(-622,11),
TO_SIGNED(-647,11),
TO_SIGNED(-670,11),
TO_SIGNED(-690,11),
TO_SIGNED(-707,11),
TO_SIGNED(-721,11),
TO_SIGNED(-733,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-731,11),
TO_SIGNED(-720,11),
TO_SIGNED(-705,11),
TO_SIGNED(-688,11),
TO_SIGNED(-667,11),
TO_SIGNED(-645,11),
TO_SIGNED(-619,11),
TO_SIGNED(-592,11),
TO_SIGNED(-562,11),
TO_SIGNED(-529,11),
TO_SIGNED(-495,11),
TO_SIGNED(-459,11),
TO_SIGNED(-421,11),
TO_SIGNED(-381,11),
TO_SIGNED(-340,11),
TO_SIGNED(-297,11),
TO_SIGNED(-254,11),
TO_SIGNED(-209,11),
TO_SIGNED(-163,11),
TO_SIGNED(-117,11),
TO_SIGNED(-70,11),
TO_SIGNED(-24,11),
TO_SIGNED(24,11),
TO_SIGNED(70,11),
TO_SIGNED(117,11),
TO_SIGNED(163,11),
TO_SIGNED(209,11),
TO_SIGNED(254,11),
TO_SIGNED(297,11),
TO_SIGNED(340,11),
TO_SIGNED(381,11),
TO_SIGNED(421,11),
TO_SIGNED(459,11),
TO_SIGNED(495,11),
TO_SIGNED(529,11),
TO_SIGNED(562,11),
TO_SIGNED(592,11),
TO_SIGNED(619,11),
TO_SIGNED(645,11),
TO_SIGNED(667,11),
TO_SIGNED(688,11),
TO_SIGNED(705,11),
TO_SIGNED(720,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(733,11),
TO_SIGNED(721,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(670,11),
TO_SIGNED(647,11),
TO_SIGNED(622,11),
TO_SIGNED(595,11),
TO_SIGNED(565,11),
TO_SIGNED(533,11),
TO_SIGNED(499,11),
TO_SIGNED(463,11),
TO_SIGNED(425,11),
TO_SIGNED(386,11),
TO_SIGNED(345,11),
TO_SIGNED(302,11),
TO_SIGNED(259,11),
TO_SIGNED(214,11),
TO_SIGNED(168,11),
TO_SIGNED(122,11),
TO_SIGNED(76,11),
TO_SIGNED(29,11),
TO_SIGNED(-18,11),
TO_SIGNED(-65,11),
TO_SIGNED(-112,11),
TO_SIGNED(-158,11),
TO_SIGNED(-204,11),
TO_SIGNED(-248,11),
TO_SIGNED(-292,11),
TO_SIGNED(-335,11),
TO_SIGNED(-376,11),
TO_SIGNED(-416,11),
TO_SIGNED(-455,11),
TO_SIGNED(-491,11),
TO_SIGNED(-526,11),
TO_SIGNED(-558,11),
TO_SIGNED(-588,11),
TO_SIGNED(-616,11),
TO_SIGNED(-642,11),
TO_SIGNED(-665,11),
TO_SIGNED(-685,11),
TO_SIGNED(-703,11),
TO_SIGNED(-718,11),
TO_SIGNED(-730,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-692,11),
TO_SIGNED(-672,11),
TO_SIGNED(-650,11),
TO_SIGNED(-625,11),
TO_SIGNED(-598,11),
TO_SIGNED(-569,11),
TO_SIGNED(-537,11),
TO_SIGNED(-503,11),
TO_SIGNED(-467,11),
TO_SIGNED(-430,11),
TO_SIGNED(-390,11),
TO_SIGNED(-349,11),
TO_SIGNED(-307,11),
TO_SIGNED(-264,11),
TO_SIGNED(-219,11),
TO_SIGNED(-174,11),
TO_SIGNED(-128,11),
TO_SIGNED(-81,11),
TO_SIGNED(-34,11),
TO_SIGNED(13,11),
TO_SIGNED(60,11),
TO_SIGNED(106,11),
TO_SIGNED(153,11),
TO_SIGNED(198,11),
TO_SIGNED(243,11),
TO_SIGNED(287,11),
TO_SIGNED(330,11),
TO_SIGNED(372,11),
TO_SIGNED(412,11),
TO_SIGNED(450,11),
TO_SIGNED(487,11),
TO_SIGNED(522,11),
TO_SIGNED(554,11),
TO_SIGNED(585,11),
TO_SIGNED(613,11),
TO_SIGNED(639,11),
TO_SIGNED(662,11),
TO_SIGNED(683,11),
TO_SIGNED(701,11),
TO_SIGNED(717,11),
TO_SIGNED(729,11),
TO_SIGNED(739,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(724,11),
TO_SIGNED(710,11),
TO_SIGNED(694,11),
TO_SIGNED(675,11),
TO_SIGNED(653,11),
TO_SIGNED(628,11),
TO_SIGNED(601,11),
TO_SIGNED(572,11),
TO_SIGNED(541,11),
TO_SIGNED(507,11),
TO_SIGNED(471,11),
TO_SIGNED(434,11),
TO_SIGNED(395,11),
TO_SIGNED(354,11),
TO_SIGNED(312,11),
TO_SIGNED(269,11),
TO_SIGNED(224,11),
TO_SIGNED(179,11),
TO_SIGNED(133,11),
TO_SIGNED(86,11),
TO_SIGNED(40,11),
TO_SIGNED(-7,11),
TO_SIGNED(-54,11),
TO_SIGNED(-101,11),
TO_SIGNED(-148,11),
TO_SIGNED(-193,11),
TO_SIGNED(-238,11),
TO_SIGNED(-282,11),
TO_SIGNED(-325,11),
TO_SIGNED(-367,11),
TO_SIGNED(-407,11),
TO_SIGNED(-446,11),
TO_SIGNED(-483,11),
TO_SIGNED(-518,11),
TO_SIGNED(-551,11),
TO_SIGNED(-582,11),
TO_SIGNED(-610,11),
TO_SIGNED(-636,11),
TO_SIGNED(-660,11),
TO_SIGNED(-681,11),
TO_SIGNED(-699,11),
TO_SIGNED(-715,11),
TO_SIGNED(-728,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-736,11),
TO_SIGNED(-725,11),
TO_SIGNED(-712,11),
TO_SIGNED(-696,11),
TO_SIGNED(-677,11),
TO_SIGNED(-655,11),
TO_SIGNED(-631,11),
TO_SIGNED(-605,11),
TO_SIGNED(-576,11),
TO_SIGNED(-544,11),
TO_SIGNED(-511,11),
TO_SIGNED(-476,11),
TO_SIGNED(-438,11),
TO_SIGNED(-399,11),
TO_SIGNED(-359,11),
TO_SIGNED(-317,11),
TO_SIGNED(-274,11),
TO_SIGNED(-229,11),
TO_SIGNED(-184,11),
TO_SIGNED(-138,11),
TO_SIGNED(-92,11),
TO_SIGNED(-45,11),
TO_SIGNED(2,11),
TO_SIGNED(49,11),
TO_SIGNED(96,11),
TO_SIGNED(142,11),
TO_SIGNED(188,11),
TO_SIGNED(233,11),
TO_SIGNED(277,11),
TO_SIGNED(321,11),
TO_SIGNED(362,11),
TO_SIGNED(403,11),
TO_SIGNED(442,11),
TO_SIGNED(479,11),
TO_SIGNED(514,11),
TO_SIGNED(547,11),
TO_SIGNED(578,11),
TO_SIGNED(607,11),
TO_SIGNED(633,11),
TO_SIGNED(657,11),
TO_SIGNED(679,11),
TO_SIGNED(697,11),
TO_SIGNED(713,11),
TO_SIGNED(726,11),
TO_SIGNED(737,11),
TO_SIGNED(744,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(744,11),
TO_SIGNED(737,11),
TO_SIGNED(727,11),
TO_SIGNED(714,11),
TO_SIGNED(698,11),
TO_SIGNED(679,11),
TO_SIGNED(658,11),
TO_SIGNED(634,11),
TO_SIGNED(608,11),
TO_SIGNED(579,11),
TO_SIGNED(548,11),
TO_SIGNED(515,11),
TO_SIGNED(480,11),
TO_SIGNED(443,11),
TO_SIGNED(404,11),
TO_SIGNED(363,11),
TO_SIGNED(322,11),
TO_SIGNED(278,11),
TO_SIGNED(234,11),
TO_SIGNED(189,11),
TO_SIGNED(143,11),
TO_SIGNED(97,11),
TO_SIGNED(50,11),
TO_SIGNED(3,11),
TO_SIGNED(-44,11),
TO_SIGNED(-91,11),
TO_SIGNED(-137,11),
TO_SIGNED(-183,11),
TO_SIGNED(-228,11),
TO_SIGNED(-273,11),
TO_SIGNED(-316,11),
TO_SIGNED(-358,11),
TO_SIGNED(-398,11),
TO_SIGNED(-437,11),
TO_SIGNED(-475,11),
TO_SIGNED(-510,11),
TO_SIGNED(-544,11),
TO_SIGNED(-575,11),
TO_SIGNED(-604,11),
TO_SIGNED(-631,11),
TO_SIGNED(-655,11),
TO_SIGNED(-676,11),
TO_SIGNED(-695,11),
TO_SIGNED(-712,11),
TO_SIGNED(-725,11),
TO_SIGNED(-736,11),
TO_SIGNED(-743,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-745,11),
TO_SIGNED(-738,11),
TO_SIGNED(-728,11),
TO_SIGNED(-715,11),
TO_SIGNED(-700,11),
TO_SIGNED(-681,11),
TO_SIGNED(-660,11),
TO_SIGNED(-637,11),
TO_SIGNED(-611,11),
TO_SIGNED(-582,11),
TO_SIGNED(-552,11),
TO_SIGNED(-519,11),
TO_SIGNED(-484,11),
TO_SIGNED(-447,11),
TO_SIGNED(-408,11),
TO_SIGNED(-368,11),
TO_SIGNED(-326,11),
TO_SIGNED(-283,11),
TO_SIGNED(-239,11),
TO_SIGNED(-194,11),
TO_SIGNED(-149,11),
TO_SIGNED(-102,11),
TO_SIGNED(-56,11),
TO_SIGNED(-9,11),
TO_SIGNED(38,11),
TO_SIGNED(85,11),
TO_SIGNED(132,11),
TO_SIGNED(178,11),
TO_SIGNED(223,11),
TO_SIGNED(268,11),
TO_SIGNED(311,11),
TO_SIGNED(353,11),
TO_SIGNED(394,11),
TO_SIGNED(433,11),
TO_SIGNED(471,11),
TO_SIGNED(506,11),
TO_SIGNED(540,11),
TO_SIGNED(571,11),
TO_SIGNED(601,11),
TO_SIGNED(628,11),
TO_SIGNED(652,11),
TO_SIGNED(674,11),
TO_SIGNED(693,11),
TO_SIGNED(710,11),
TO_SIGNED(724,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(739,11),
TO_SIGNED(729,11),
TO_SIGNED(717,11),
TO_SIGNED(702,11),
TO_SIGNED(684,11),
TO_SIGNED(663,11),
TO_SIGNED(640,11),
TO_SIGNED(614,11),
TO_SIGNED(586,11),
TO_SIGNED(555,11),
TO_SIGNED(523,11),
TO_SIGNED(488,11),
TO_SIGNED(451,11),
TO_SIGNED(413,11),
TO_SIGNED(373,11),
TO_SIGNED(331,11),
TO_SIGNED(288,11),
TO_SIGNED(244,11),
TO_SIGNED(200,11),
TO_SIGNED(154,11),
TO_SIGNED(108,11),
TO_SIGNED(61,11),
TO_SIGNED(14,11),
TO_SIGNED(-33,11),
TO_SIGNED(-80,11),
TO_SIGNED(-127,11),
TO_SIGNED(-173,11),
TO_SIGNED(-218,11),
TO_SIGNED(-263,11),
TO_SIGNED(-306,11),
TO_SIGNED(-348,11),
TO_SIGNED(-389,11),
TO_SIGNED(-429,11),
TO_SIGNED(-466,11),
TO_SIGNED(-502,11),
TO_SIGNED(-536,11),
TO_SIGNED(-568,11),
TO_SIGNED(-598,11),
TO_SIGNED(-625,11),
TO_SIGNED(-650,11),
TO_SIGNED(-672,11),
TO_SIGNED(-691,11),
TO_SIGNED(-708,11),
TO_SIGNED(-722,11),
TO_SIGNED(-733,11),
TO_SIGNED(-742,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-740,11),
TO_SIGNED(-730,11),
TO_SIGNED(-718,11),
TO_SIGNED(-703,11),
TO_SIGNED(-686,11),
TO_SIGNED(-665,11),
TO_SIGNED(-642,11),
TO_SIGNED(-617,11),
TO_SIGNED(-589,11),
TO_SIGNED(-559,11),
TO_SIGNED(-526,11),
TO_SIGNED(-492,11),
TO_SIGNED(-455,11),
TO_SIGNED(-417,11),
TO_SIGNED(-377,11),
TO_SIGNED(-336,11),
TO_SIGNED(-293,11),
TO_SIGNED(-249,11),
TO_SIGNED(-205,11),
TO_SIGNED(-159,11),
TO_SIGNED(-113,11),
TO_SIGNED(-66,11),
TO_SIGNED(-19,11),
TO_SIGNED(28,11),
TO_SIGNED(75,11),
TO_SIGNED(121,11),
TO_SIGNED(167,11),
TO_SIGNED(213,11),
TO_SIGNED(258,11),
TO_SIGNED(301,11),
TO_SIGNED(344,11),
TO_SIGNED(385,11),
TO_SIGNED(424,11),
TO_SIGNED(462,11),
TO_SIGNED(498,11),
TO_SIGNED(532,11),
TO_SIGNED(564,11),
TO_SIGNED(594,11),
TO_SIGNED(622,11),
TO_SIGNED(647,11),
TO_SIGNED(669,11),
TO_SIGNED(689,11),
TO_SIGNED(706,11),
TO_SIGNED(721,11),
TO_SIGNED(732,11),
TO_SIGNED(741,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(741,11),
TO_SIGNED(732,11),
TO_SIGNED(720,11),
TO_SIGNED(705,11),
TO_SIGNED(688,11),
TO_SIGNED(668,11),
TO_SIGNED(645,11),
TO_SIGNED(620,11),
TO_SIGNED(592,11),
TO_SIGNED(562,11),
TO_SIGNED(530,11),
TO_SIGNED(496,11),
TO_SIGNED(460,11),
TO_SIGNED(422,11),
TO_SIGNED(382,11),
TO_SIGNED(341,11),
TO_SIGNED(298,11),
TO_SIGNED(255,11),
TO_SIGNED(210,11),
TO_SIGNED(164,11),
TO_SIGNED(118,11),
TO_SIGNED(71,11),
TO_SIGNED(25,11),
TO_SIGNED(-22,11),
TO_SIGNED(-69,11),
TO_SIGNED(-116,11),
TO_SIGNED(-162,11),
TO_SIGNED(-208,11),
TO_SIGNED(-252,11),
TO_SIGNED(-296,11),
TO_SIGNED(-339,11),
TO_SIGNED(-380,11),
TO_SIGNED(-420,11),
TO_SIGNED(-458,11),
TO_SIGNED(-494,11),
TO_SIGNED(-529,11),
TO_SIGNED(-561,11),
TO_SIGNED(-591,11),
TO_SIGNED(-619,11),
TO_SIGNED(-644,11),
TO_SIGNED(-667,11),
TO_SIGNED(-687,11),
TO_SIGNED(-705,11),
TO_SIGNED(-719,11),
TO_SIGNED(-731,11),
TO_SIGNED(-740,11),
TO_SIGNED(-746,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-733,11),
TO_SIGNED(-721,11),
TO_SIGNED(-707,11),
TO_SIGNED(-690,11),
TO_SIGNED(-670,11),
TO_SIGNED(-648,11),
TO_SIGNED(-623,11),
TO_SIGNED(-596,11),
TO_SIGNED(-566,11),
TO_SIGNED(-534,11),
TO_SIGNED(-500,11),
TO_SIGNED(-464,11),
TO_SIGNED(-426,11),
TO_SIGNED(-387,11),
TO_SIGNED(-345,11),
TO_SIGNED(-303,11),
TO_SIGNED(-260,11),
TO_SIGNED(-215,11),
TO_SIGNED(-169,11),
TO_SIGNED(-123,11),
TO_SIGNED(-77,11),
TO_SIGNED(-30,11),
TO_SIGNED(17,11),
TO_SIGNED(64,11),
TO_SIGNED(111,11),
TO_SIGNED(157,11),
TO_SIGNED(203,11),
TO_SIGNED(247,11),
TO_SIGNED(291,11),
TO_SIGNED(334,11),
TO_SIGNED(375,11),
TO_SIGNED(415,11),
TO_SIGNED(454,11),
TO_SIGNED(490,11),
TO_SIGNED(525,11),
TO_SIGNED(557,11),
TO_SIGNED(588,11),
TO_SIGNED(616,11),
TO_SIGNED(641,11),
TO_SIGNED(664,11),
TO_SIGNED(685,11),
TO_SIGNED(703,11),
TO_SIGNED(718,11),
TO_SIGNED(730,11),
TO_SIGNED(739,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(734,11),
TO_SIGNED(723,11),
TO_SIGNED(709,11),
TO_SIGNED(692,11),
TO_SIGNED(673,11),
TO_SIGNED(651,11),
TO_SIGNED(626,11),
TO_SIGNED(599,11),
TO_SIGNED(569,11),
TO_SIGNED(538,11),
TO_SIGNED(504,11),
TO_SIGNED(468,11),
TO_SIGNED(430,11),
TO_SIGNED(391,11),
TO_SIGNED(350,11),
TO_SIGNED(308,11),
TO_SIGNED(265,11),
TO_SIGNED(220,11),
TO_SIGNED(175,11),
TO_SIGNED(129,11),
TO_SIGNED(82,11),
TO_SIGNED(35,11),
TO_SIGNED(-12,11),
TO_SIGNED(-59,11),
TO_SIGNED(-105,11),
TO_SIGNED(-152,11),
TO_SIGNED(-197,11),
TO_SIGNED(-242,11),
TO_SIGNED(-286,11),
TO_SIGNED(-329,11),
TO_SIGNED(-371,11),
TO_SIGNED(-411,11),
TO_SIGNED(-449,11),
TO_SIGNED(-486,11),
TO_SIGNED(-521,11),
TO_SIGNED(-554,11),
TO_SIGNED(-584,11),
TO_SIGNED(-613,11),
TO_SIGNED(-639,11),
TO_SIGNED(-662,11),
TO_SIGNED(-683,11),
TO_SIGNED(-701,11),
TO_SIGNED(-716,11),
TO_SIGNED(-729,11),
TO_SIGNED(-738,11),
TO_SIGNED(-745,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-743,11),
TO_SIGNED(-735,11),
TO_SIGNED(-724,11),
TO_SIGNED(-711,11),
TO_SIGNED(-694,11),
TO_SIGNED(-675,11),
TO_SIGNED(-653,11),
TO_SIGNED(-629,11),
TO_SIGNED(-602,11),
TO_SIGNED(-573,11),
TO_SIGNED(-541,11),
TO_SIGNED(-508,11),
TO_SIGNED(-472,11),
TO_SIGNED(-435,11),
TO_SIGNED(-396,11),
TO_SIGNED(-355,11),
TO_SIGNED(-313,11),
TO_SIGNED(-270,11),
TO_SIGNED(-225,11),
TO_SIGNED(-180,11),
TO_SIGNED(-134,11),
TO_SIGNED(-87,11),
TO_SIGNED(-41,11),
TO_SIGNED(6,11),
TO_SIGNED(53,11),
TO_SIGNED(100,11),
TO_SIGNED(147,11),
TO_SIGNED(192,11),
TO_SIGNED(237,11),
TO_SIGNED(281,11),
TO_SIGNED(324,11),
TO_SIGNED(366,11),
TO_SIGNED(406,11),
TO_SIGNED(445,11),
TO_SIGNED(482,11),
TO_SIGNED(517,11),
TO_SIGNED(550,11),
TO_SIGNED(581,11),
TO_SIGNED(610,11),
TO_SIGNED(636,11),
TO_SIGNED(659,11),
TO_SIGNED(681,11),
TO_SIGNED(699,11),
TO_SIGNED(715,11),
TO_SIGNED(727,11),
TO_SIGNED(737,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(744,11),
TO_SIGNED(736,11),
TO_SIGNED(726,11),
TO_SIGNED(712,11),
TO_SIGNED(696,11),
TO_SIGNED(677,11),
TO_SIGNED(656,11),
TO_SIGNED(632,11),
TO_SIGNED(605,11),
TO_SIGNED(576,11),
TO_SIGNED(545,11),
TO_SIGNED(512,11),
TO_SIGNED(476,11),
TO_SIGNED(439,11),
TO_SIGNED(400,11),
TO_SIGNED(360,11),
TO_SIGNED(318,11),
TO_SIGNED(275,11),
TO_SIGNED(230,11),
TO_SIGNED(185,11),
TO_SIGNED(139,11),
TO_SIGNED(93,11),
TO_SIGNED(46,11),
TO_SIGNED(-1,11),
TO_SIGNED(-48,11),
TO_SIGNED(-95,11),
TO_SIGNED(-141,11),
TO_SIGNED(-187,11),
TO_SIGNED(-232,11),
TO_SIGNED(-276,11),
TO_SIGNED(-320,11),
TO_SIGNED(-362,11),
TO_SIGNED(-402,11),
TO_SIGNED(-441,11),
TO_SIGNED(-478,11),
TO_SIGNED(-513,11),
TO_SIGNED(-547,11),
TO_SIGNED(-578,11),
TO_SIGNED(-606,11),
TO_SIGNED(-633,11),
TO_SIGNED(-657,11),
TO_SIGNED(-678,11),
TO_SIGNED(-697,11),
TO_SIGNED(-713,11),
TO_SIGNED(-726,11),
TO_SIGNED(-736,11),
TO_SIGNED(-744,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-744,11),
TO_SIGNED(-737,11),
TO_SIGNED(-727,11),
TO_SIGNED(-714,11),
TO_SIGNED(-698,11),
TO_SIGNED(-680,11),
TO_SIGNED(-658,11),
TO_SIGNED(-635,11),
TO_SIGNED(-608,11),
TO_SIGNED(-580,11),
TO_SIGNED(-549,11),
TO_SIGNED(-516,11),
TO_SIGNED(-480,11),
TO_SIGNED(-443,11),
TO_SIGNED(-405,11),
TO_SIGNED(-364,11),
TO_SIGNED(-323,11),
TO_SIGNED(-279,11),
TO_SIGNED(-235,11),
TO_SIGNED(-190,11),
TO_SIGNED(-144,11),
TO_SIGNED(-98,11),
TO_SIGNED(-51,11),
TO_SIGNED(-4,11),
TO_SIGNED(43,11),
TO_SIGNED(90,11),
TO_SIGNED(136,11),
TO_SIGNED(182,11),
TO_SIGNED(227,11),
TO_SIGNED(272,11),
TO_SIGNED(315,11),
TO_SIGNED(357,11),
TO_SIGNED(397,11),
TO_SIGNED(437,11),
TO_SIGNED(474,11),
TO_SIGNED(509,11),
TO_SIGNED(543,11),
TO_SIGNED(574,11),
TO_SIGNED(603,11),
TO_SIGNED(630,11),
TO_SIGNED(654,11),
TO_SIGNED(676,11),
TO_SIGNED(695,11),
TO_SIGNED(711,11),
TO_SIGNED(725,11),
TO_SIGNED(735,11),
TO_SIGNED(743,11),
TO_SIGNED(748,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(745,11),
TO_SIGNED(738,11),
TO_SIGNED(728,11),
TO_SIGNED(716,11),
TO_SIGNED(700,11),
TO_SIGNED(682,11),
TO_SIGNED(661,11),
TO_SIGNED(637,11),
TO_SIGNED(611,11),
TO_SIGNED(583,11),
TO_SIGNED(552,11),
TO_SIGNED(519,11),
TO_SIGNED(485,11),
TO_SIGNED(448,11),
TO_SIGNED(409,11),
TO_SIGNED(369,11),
TO_SIGNED(327,11),
TO_SIGNED(284,11),
TO_SIGNED(240,11),
TO_SIGNED(195,11),
TO_SIGNED(150,11),
TO_SIGNED(103,11),
TO_SIGNED(57,11),
TO_SIGNED(10,11),
TO_SIGNED(-37,11),
TO_SIGNED(-84,11),
TO_SIGNED(-131,11),
TO_SIGNED(-177,11),
TO_SIGNED(-222,11),
TO_SIGNED(-267,11),
TO_SIGNED(-310,11),
TO_SIGNED(-352,11),
TO_SIGNED(-393,11),
TO_SIGNED(-432,11),
TO_SIGNED(-470,11),
TO_SIGNED(-505,11),
TO_SIGNED(-539,11),
TO_SIGNED(-571,11),
TO_SIGNED(-600,11),
TO_SIGNED(-627,11),
TO_SIGNED(-652,11),
TO_SIGNED(-674,11),
TO_SIGNED(-693,11),
TO_SIGNED(-710,11),
TO_SIGNED(-723,11),
TO_SIGNED(-734,11),
TO_SIGNED(-742,11),
TO_SIGNED(-748,11),
TO_SIGNED(-750,11),
TO_SIGNED(-749,11),
TO_SIGNED(-746,11),
TO_SIGNED(-739,11),
TO_SIGNED(-729,11),
TO_SIGNED(-717,11),
TO_SIGNED(-702,11),
TO_SIGNED(-684,11),
TO_SIGNED(-663,11),
TO_SIGNED(-640,11),
TO_SIGNED(-615,11),
TO_SIGNED(-586,11),
TO_SIGNED(-556,11),
TO_SIGNED(-523,11),
TO_SIGNED(-489,11),
TO_SIGNED(-452,11),
TO_SIGNED(-414,11),
TO_SIGNED(-374,11),
TO_SIGNED(-332,11),
TO_SIGNED(-289,11),
TO_SIGNED(-245,11),
TO_SIGNED(-201,11),
TO_SIGNED(-155,11),
TO_SIGNED(-109,11),
TO_SIGNED(-62,11),
TO_SIGNED(-15,11),
TO_SIGNED(32,11),
TO_SIGNED(79,11),
TO_SIGNED(125,11),
TO_SIGNED(172,11),
TO_SIGNED(217,11),
TO_SIGNED(262,11),
TO_SIGNED(305,11),
TO_SIGNED(347,11),
TO_SIGNED(388,11),
TO_SIGNED(428,11),
TO_SIGNED(466,11),
TO_SIGNED(501,11),
TO_SIGNED(535,11),
TO_SIGNED(567,11),
TO_SIGNED(597,11),
TO_SIGNED(624,11),
TO_SIGNED(649,11),
TO_SIGNED(671,11),
TO_SIGNED(691,11),
TO_SIGNED(708,11),
TO_SIGNED(722,11),
TO_SIGNED(733,11),
TO_SIGNED(742,11),
TO_SIGNED(747,11),
TO_SIGNED(750,11),
TO_SIGNED(749,11),
TO_SIGNED(746,11),
TO_SIGNED(740,11),
TO_SIGNED(731,11),
TO_SIGNED(719,11),
TO_SIGNED(704,11),
TO_SIGNED(686,11),
TO_SIGNED(666,11),
TO_SIGNED(643,11),
TO_SIGNED(618,11),
TO_SIGNED(590,11),
TO_SIGNED(559,11),
TO_SIGNED(527,11),
TO_SIGNED(493,11),
TO_SIGNED(456,11),
TO_SIGNED(418,11),
TO_SIGNED(378,11),
TO_SIGNED(337,11),
TO_SIGNED(294,11),
TO_SIGNED(250,11),
TO_SIGNED(206,11),
TO_SIGNED(160,11),
TO_SIGNED(114,11),
TO_SIGNED(67,11),
TO_SIGNED(20,11),
TO_SIGNED(-27,11),
TO_SIGNED(-74,11),
TO_SIGNED(-120,11),
TO_SIGNED(-166,11),
TO_SIGNED(-212,11),
TO_SIGNED(-257,11),
TO_SIGNED(-300,11),
TO_SIGNED(-343,11),
TO_SIGNED(-384,11),
TO_SIGNED(-423,11),
TO_SIGNED(-461,11),
TO_SIGNED(-497,11),
TO_SIGNED(-532,11),
TO_SIGNED(-564,11),
TO_SIGNED(-594,11),
TO_SIGNED(-621,11),
TO_SIGNED(-646,11),
TO_SIGNED(-669,11),
TO_SIGNED(-689,11),
TO_SIGNED(-706,11),
TO_SIGNED(-721,11),
TO_SIGNED(-732,11),
TO_SIGNED(-741,11),
TO_SIGNED(-747,11),
TO_SIGNED(-750,11),
TO_SIGNED(-750,11),
TO_SIGNED(-747,11),
TO_SIGNED(-741,11),
TO_SIGNED(-732,11),
TO_SIGNED(-720,11),
TO_SIGNED(-706,11),
TO_SIGNED(-688,11),
TO_SIGNED(-668,11),
TO_SIGNED(-646,11),
TO_SIGNED(-621,11),
TO_SIGNED(-593,11),
TO_SIGNED(-563,11),
TO_SIGNED(-531,11),
TO_SIGNED(-497,11),
TO_SIGNED(-460,11),
TO_SIGNED(-422,11),
TO_SIGNED(-383,11),
TO_SIGNED(-342,11),
TO_SIGNED(-299,11),
TO_SIGNED(-256,11),
TO_SIGNED(-211,11),
TO_SIGNED(-165,11),
TO_SIGNED(-119,11),
TO_SIGNED(-73,11),
TO_SIGNED(-26,11),
TO_SIGNED(21,11),
TO_SIGNED(68,11),
TO_SIGNED(115,11),
TO_SIGNED(161,11),
TO_SIGNED(207,11),
TO_SIGNED(251,11),
TO_SIGNED(295,11),
TO_SIGNED(338,11),
TO_SIGNED(379,11),
TO_SIGNED(419,11),
TO_SIGNED(457,11),
TO_SIGNED(493,11),
TO_SIGNED(528,11),
TO_SIGNED(560,11),
TO_SIGNED(590,11),
TO_SIGNED(618,11),
TO_SIGNED(644,11),
TO_SIGNED(666,11),
TO_SIGNED(687,11),
TO_SIGNED(704,11),
TO_SIGNED(719,11),
TO_SIGNED(731,11),
TO_SIGNED(740,11),
TO_SIGNED(746,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(747,11),
TO_SIGNED(742,11),
TO_SIGNED(733,11),
TO_SIGNED(722,11),
TO_SIGNED(707,11),
TO_SIGNED(690,11),
TO_SIGNED(671,11),
TO_SIGNED(648,11),
TO_SIGNED(624,11),
TO_SIGNED(596,11),
TO_SIGNED(567,11),
TO_SIGNED(535,11),
TO_SIGNED(501,11),
TO_SIGNED(465,11),
TO_SIGNED(427,11),
TO_SIGNED(387,11),
TO_SIGNED(346,11),
TO_SIGNED(304,11),
TO_SIGNED(261,11),
TO_SIGNED(216,11),
TO_SIGNED(171,11),
TO_SIGNED(124,11),
TO_SIGNED(78,11),
TO_SIGNED(31,11),
TO_SIGNED(-16,11),
TO_SIGNED(-63,11),
TO_SIGNED(-110,11),
TO_SIGNED(-156,11),
TO_SIGNED(-202,11),
TO_SIGNED(-246,11),
TO_SIGNED(-290,11),
TO_SIGNED(-333,11),
TO_SIGNED(-375,11),
TO_SIGNED(-415,11),
TO_SIGNED(-453,11),
TO_SIGNED(-489,11),
TO_SIGNED(-524,11),
TO_SIGNED(-557,11),
TO_SIGNED(-587,11),
TO_SIGNED(-615,11),
TO_SIGNED(-641,11),
TO_SIGNED(-664,11),
TO_SIGNED(-685,11),
TO_SIGNED(-702,11),
TO_SIGNED(-717,11),
TO_SIGNED(-730,11),
TO_SIGNED(-739,11),
TO_SIGNED(-746,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-742,11),
TO_SIGNED(-734,11),
TO_SIGNED(-723,11),
TO_SIGNED(-709,11),
TO_SIGNED(-693,11),
TO_SIGNED(-673,11),
TO_SIGNED(-651,11),
TO_SIGNED(-627,11),
TO_SIGNED(-599,11),
TO_SIGNED(-570,11),
TO_SIGNED(-538,11),
TO_SIGNED(-505,11),
TO_SIGNED(-469,11),
TO_SIGNED(-431,11),
TO_SIGNED(-392,11),
TO_SIGNED(-351,11),
TO_SIGNED(-309,11),
TO_SIGNED(-266,11),
TO_SIGNED(-221,11),
TO_SIGNED(-176,11),
TO_SIGNED(-130,11),
TO_SIGNED(-83,11),
TO_SIGNED(-36,11),
TO_SIGNED(11,11),
TO_SIGNED(58,11),
TO_SIGNED(104,11),
TO_SIGNED(151,11),
TO_SIGNED(196,11),
TO_SIGNED(241,11),
TO_SIGNED(285,11),
TO_SIGNED(328,11),
TO_SIGNED(370,11),
TO_SIGNED(410,11),
TO_SIGNED(449,11),
TO_SIGNED(485,11),
TO_SIGNED(520,11),
TO_SIGNED(553,11),
TO_SIGNED(584,11),
TO_SIGNED(612,11),
TO_SIGNED(638,11),
TO_SIGNED(661,11),
TO_SIGNED(682,11),
TO_SIGNED(700,11),
TO_SIGNED(716,11),
TO_SIGNED(728,11),
TO_SIGNED(738,11),
TO_SIGNED(745,11),
TO_SIGNED(749,11),
TO_SIGNED(750,11),
TO_SIGNED(748,11),
TO_SIGNED(743,11),
TO_SIGNED(735,11),
TO_SIGNED(725,11),
TO_SIGNED(711,11),
TO_SIGNED(695,11),
TO_SIGNED(675,11),
TO_SIGNED(654,11),
TO_SIGNED(629,11),
TO_SIGNED(603,11),
TO_SIGNED(574,11),
TO_SIGNED(542,11),
TO_SIGNED(509,11),
TO_SIGNED(473,11),
TO_SIGNED(436,11),
TO_SIGNED(397,11),
TO_SIGNED(356,11),
TO_SIGNED(314,11),
TO_SIGNED(271,11),
TO_SIGNED(226,11),
TO_SIGNED(181,11),
TO_SIGNED(135,11),
TO_SIGNED(88,11),
TO_SIGNED(42,11),
TO_SIGNED(-5,11),
TO_SIGNED(-52,11),
TO_SIGNED(-99,11),
TO_SIGNED(-145,11),
TO_SIGNED(-191,11),
TO_SIGNED(-236,11),
TO_SIGNED(-280,11),
TO_SIGNED(-323,11),
TO_SIGNED(-365,11),
TO_SIGNED(-406,11),
TO_SIGNED(-444,11),
TO_SIGNED(-481,11),
TO_SIGNED(-516,11),
TO_SIGNED(-549,11),
TO_SIGNED(-580,11),
TO_SIGNED(-609,11),
TO_SIGNED(-635,11),
TO_SIGNED(-659,11),
TO_SIGNED(-680,11),
TO_SIGNED(-699,11),
TO_SIGNED(-714,11),
TO_SIGNED(-727,11),
TO_SIGNED(-737,11),
TO_SIGNED(-744,11),
TO_SIGNED(-749,11),
TO_SIGNED(-750,11),
TO_SIGNED(-748,11),
TO_SIGNED(-744,11),
TO_SIGNED(-736,11),
TO_SIGNED(-726,11),
TO_SIGNED(-713,11),
TO_SIGNED(-697,11),
TO_SIGNED(-678,11),
TO_SIGNED(-656,11),
TO_SIGNED(-632,11),
TO_SIGNED(-606,11),
TO_SIGNED(-577,11),
TO_SIGNED(-546,11),
TO_SIGNED(-512,11),
TO_SIGNED(-477,11),
TO_SIGNED(-440,11),
TO_SIGNED(-401,11),
TO_SIGNED(-361,11),
TO_SIGNED(-319,11),
TO_SIGNED(-275,11),
TO_SIGNED(-231,11),
TO_SIGNED(-186,11),
TO_SIGNED(-140,11),
TO_SIGNED(-94,11),
TO_SIGNED(-47,11)
  );

signal data_n1, data_n2 : std_logic_vector(10 downto 0);
signal sum_div2 : unsigned(10 downto 0);

BEGIN
PROCESS (CLOCK)
BEGIN
IF RISING_EDGE(CLOCK) THEN
    if(ce  = '1') then
    
    data_n1 <= STD_LOGIC_VECTOR(memory(TO_INTEGER(unsigned(addr_1))));
    IF two_notes = '1' THEN
        data_n2 <= STD_LOGIC_VECTOR(memory(TO_INTEGER(unsigned(addr_2))));
    ELSE
        data_n2 <= (others => '0'); 
    END IF;

  
    IF two_notes = '1' THEN
       
        sum_div2 <= (unsigned(data_n1) + unsigned(data_n2)) srl 1; 
        DATA_OUT <=std_logic_vector(sum_div2);
    ELSE
        
        DATA_OUT <= data_n1;
    END IF;
END IF;
end if;
END PROCESS;



END Behavioral;